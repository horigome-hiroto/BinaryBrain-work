`timescale 1ns / 1ps



module MnistLutSimple
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire                  reset,
            input  wire                  clk,
            input  wire                  cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [      784-1:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [       10-1:0]  out_data,
            output wire                  out_valid
        );
    
    
    wire  [USER_BITS-1:0]  layer0_user;
    wire  [     2304-1:0]  layer0_data;
    wire                   layer0_valid;
    
    MnistLutSimple_sub0
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub0
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (in_user),
                .in_data    (in_data),
                .in_valid   (in_valid),
                
                .out_user   (layer0_user),
                .out_data   (layer0_data),
                .out_valid  (layer0_valid)
             );
    
    wire  [USER_BITS-1:0]  layer1_user;
    wire  [      384-1:0]  layer1_data;
    wire                   layer1_valid;
    
    MnistLutSimple_sub1
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub1
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer0_user),
                .in_data    (layer0_data),
                .in_valid   (layer0_valid),
                
                .out_user   (layer1_user),
                .out_data   (layer1_data),
                .out_valid  (layer1_valid)
             );
    
    wire  [USER_BITS-1:0]  layer2_user;
    wire  [       64-1:0]  layer2_data;
    wire                   layer2_valid;
    
    MnistLutSimple_sub2
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub2
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer1_user),
                .in_data    (layer1_data),
                .in_valid   (layer1_valid),
                
                .out_user   (layer2_user),
                .out_data   (layer2_data),
                .out_valid  (layer2_valid)
             );
    
    wire  [USER_BITS-1:0]  layer3_user;
    wire  [      360-1:0]  layer3_data;
    wire                   layer3_valid;
    
    MnistLutSimple_sub3
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub3
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer2_user),
                .in_data    (layer2_data),
                .in_valid   (layer2_valid),
                
                .out_user   (layer3_user),
                .out_data   (layer3_data),
                .out_valid  (layer3_valid)
             );
    
    wire  [USER_BITS-1:0]  layer4_user;
    wire  [       60-1:0]  layer4_data;
    wire                   layer4_valid;
    
    MnistLutSimple_sub4
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub4
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer3_user),
                .in_data    (layer3_data),
                .in_valid   (layer3_valid),
                
                .out_user   (layer4_user),
                .out_data   (layer4_data),
                .out_valid  (layer4_valid)
             );
    
    wire  [USER_BITS-1:0]  layer5_user;
    wire  [       10-1:0]  layer5_data;
    wire                   layer5_valid;
    
    MnistLutSimple_sub5
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub5
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer4_user),
                .in_data    (layer4_data),
                .in_valid   (layer4_valid),
                
                .out_user   (layer5_user),
                .out_data   (layer5_data),
                .out_valid  (layer5_valid)
             );
    
    assign out_data  = layer5_data;
    assign out_user  = layer5_user;
    assign out_valid = layer5_valid;
    
endmodule




module MnistLutSimple_sub0
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        783:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [       2303:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub0_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub0_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub0_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [783:0]  in_data,
            output wire [2303:0]  out_data
        );
    
    
    // LUT : 0
    wire [63:0] lut_0_table = 64'b1111110011111100111111001101110011111100111111001101110011011100;
    wire [5:0] lut_0_select = {
                             in_data[111],
                             in_data[736],
                             in_data[420],
                             in_data[316],
                             in_data[302],
                             in_data[531]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [63:0] lut_1_table = 64'b1100111101001111000000000100110011001111010011110000100001001100;
    wire [5:0] lut_1_select = {
                             in_data[20],
                             in_data[400],
                             in_data[203],
                             in_data[529],
                             in_data[191],
                             in_data[73]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [63:0] lut_2_table = 64'b1111111111111111100011111000111011111111111111111010111010101110;
    wire [5:0] lut_2_select = {
                             in_data[310],
                             in_data[148],
                             in_data[725],
                             in_data[692],
                             in_data[677],
                             in_data[620]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [63:0] lut_3_table = 64'b0000000010101010101010101111101100000000111111111010100011111010;
    wire [5:0] lut_3_select = {
                             in_data[330],
                             in_data[606],
                             in_data[98],
                             in_data[501],
                             in_data[44],
                             in_data[663]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [63:0] lut_4_table = 64'b1111111111111111111111001111111111111111111111111100110011111111;
    wire [5:0] lut_4_select = {
                             in_data[132],
                             in_data[707],
                             in_data[428],
                             in_data[129],
                             in_data[742],
                             in_data[334]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [63:0] lut_5_table = 64'b0011010111111101001101010111110100110011001100110011001100110011;
    wire [5:0] lut_5_select = {
                             in_data[574],
                             in_data[419],
                             in_data[699],
                             in_data[193],
                             in_data[298],
                             in_data[771]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [63:0] lut_6_table = 64'b0000000011000000110000001100110000000000110011001100110111111111;
    wire [5:0] lut_6_select = {
                             in_data[414],
                             in_data[359],
                             in_data[580],
                             in_data[40],
                             in_data[608],
                             in_data[783]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [63:0] lut_7_table = 64'b1111111111111111010011001100110011111111111111111100110011001100;
    wire [5:0] lut_7_select = {
                             in_data[338],
                             in_data[397],
                             in_data[424],
                             in_data[502],
                             in_data[320],
                             in_data[696]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [63:0] lut_8_table = 64'b0000000011110101000001011101010110000000111101010000010111010101;
    wire [5:0] lut_8_select = {
                             in_data[394],
                             in_data[101],
                             in_data[512],
                             in_data[490],
                             in_data[480],
                             in_data[433]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [63:0] lut_9_table = 64'b1010101000001010000011110000111010101010000010101111111100001111;
    wire [5:0] lut_9_select = {
                             in_data[585],
                             in_data[322],
                             in_data[745],
                             in_data[472],
                             in_data[141],
                             in_data[355]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [63:0] lut_10_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_10_select = {
                             in_data[561],
                             in_data[629],
                             in_data[252],
                             in_data[522],
                             in_data[753],
                             in_data[296]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [63:0] lut_11_table = 64'b0000000000000000000000000000000000000100111111110101010101010101;
    wire [5:0] lut_11_select = {
                             in_data[125],
                             in_data[426],
                             in_data[483],
                             in_data[560],
                             in_data[53],
                             in_data[689]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [63:0] lut_12_table = 64'b1111111111111111000011010000111101000101010011010000010100001101;
    wire [5:0] lut_12_select = {
                             in_data[123],
                             in_data[147],
                             in_data[340],
                             in_data[602],
                             in_data[171],
                             in_data[470]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [63:0] lut_13_table = 64'b0011001100110001000000010000000011111111111111110001010100010001;
    wire [5:0] lut_13_select = {
                             in_data[513],
                             in_data[690],
                             in_data[767],
                             in_data[168],
                             in_data[128],
                             in_data[232]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [63:0] lut_14_table = 64'b0000000001011111000000000000010111011111111111110000000001011111;
    wire [5:0] lut_14_select = {
                             in_data[526],
                             in_data[276],
                             in_data[352],
                             in_data[104],
                             in_data[19],
                             in_data[94]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [63:0] lut_15_table = 64'b1111111101000000111111111100000011111111110001001111111111001100;
    wire [5:0] lut_15_select = {
                             in_data[600],
                             in_data[79],
                             in_data[267],
                             in_data[485],
                             in_data[446],
                             in_data[701]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [63:0] lut_16_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_16_select = {
                             in_data[353],
                             in_data[116],
                             in_data[337],
                             in_data[58],
                             in_data[97],
                             in_data[368]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [63:0] lut_17_table = 64'b1111111111111111111110111111111110110000101100101111001011110010;
    wire [5:0] lut_17_select = {
                             in_data[304],
                             in_data[221],
                             in_data[738],
                             in_data[481],
                             in_data[749],
                             in_data[77]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [63:0] lut_18_table = 64'b0111011101110111111111111111111100000000000000000101110111010101;
    wire [5:0] lut_18_select = {
                             in_data[152],
                             in_data[216],
                             in_data[33],
                             in_data[167],
                             in_data[374],
                             in_data[506]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [63:0] lut_19_table = 64'b0000000000000000000000000000000000000000111111110000000011111111;
    wire [5:0] lut_19_select = {
                             in_data[605],
                             in_data[389],
                             in_data[565],
                             in_data[728],
                             in_data[365],
                             in_data[166]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [63:0] lut_20_table = 64'b0010000011110000111100001111001100110000111100001111000011110011;
    wire [5:0] lut_20_select = {
                             in_data[64],
                             in_data[545],
                             in_data[436],
                             in_data[427],
                             in_data[172],
                             in_data[393]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [63:0] lut_21_table = 64'b0000000010101111101010101010111100000000101011111010101010101111;
    wire [5:0] lut_21_select = {
                             in_data[54],
                             in_data[435],
                             in_data[549],
                             in_data[662],
                             in_data[26],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [63:0] lut_22_table = 64'b0000000000110101000000000001000100000000001101010000000000110001;
    wire [5:0] lut_22_select = {
                             in_data[43],
                             in_data[107],
                             in_data[444],
                             in_data[628],
                             in_data[332],
                             in_data[431]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [63:0] lut_23_table = 64'b1100110011001100000011001100110011001100110011001100110011001100;
    wire [5:0] lut_23_select = {
                             in_data[648],
                             in_data[719],
                             in_data[195],
                             in_data[622],
                             in_data[489],
                             in_data[35]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [63:0] lut_24_table = 64'b1111111111111111111111111011101111111111001100111011101110100000;
    wire [5:0] lut_24_select = {
                             in_data[511],
                             in_data[155],
                             in_data[510],
                             in_data[724],
                             in_data[403],
                             in_data[269]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [63:0] lut_25_table = 64'b0000000000000000101010101011101100000000000000001010101010101010;
    wire [5:0] lut_25_select = {
                             in_data[63],
                             in_data[459],
                             in_data[504],
                             in_data[142],
                             in_data[176],
                             in_data[601]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [63:0] lut_26_table = 64'b1100110011111111000100001111111111001100110011100000000011111111;
    wire [5:0] lut_26_select = {
                             in_data[361],
                             in_data[236],
                             in_data[434],
                             in_data[718],
                             in_data[179],
                             in_data[131]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [63:0] lut_27_table = 64'b1101110100000100110011000000000011111111100011011100110000000000;
    wire [5:0] lut_27_select = {
                             in_data[717],
                             in_data[164],
                             in_data[494],
                             in_data[223],
                             in_data[521],
                             in_data[432]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [63:0] lut_28_table = 64'b0000000000000000000000000000000000000101000001010000010100000101;
    wire [5:0] lut_28_select = {
                             in_data[678],
                             in_data[774],
                             in_data[84],
                             in_data[634],
                             in_data[2],
                             in_data[528]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [63:0] lut_29_table = 64'b0000111100001111000001110000000000001111000011110000111100001111;
    wire [5:0] lut_29_select = {
                             in_data[706],
                             in_data[130],
                             in_data[186],
                             in_data[488],
                             in_data[42],
                             in_data[331]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [63:0] lut_30_table = 64'b0000000011001100000000001100000011111100111111011111100011111100;
    wire [5:0] lut_30_select = {
                             in_data[286],
                             in_data[99],
                             in_data[415],
                             in_data[333],
                             in_data[151],
                             in_data[576]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [63:0] lut_31_table = 64'b0000000000000000000000010000000000000000000000001111111100001111;
    wire [5:0] lut_31_select = {
                             in_data[228],
                             in_data[408],
                             in_data[160],
                             in_data[437],
                             in_data[779],
                             in_data[649]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [63:0] lut_32_table = 64'b0000000000110000000000001111000000000000001100000000000011110000;
    wire [5:0] lut_32_select = {
                             in_data[60],
                             in_data[465],
                             in_data[294],
                             in_data[402],
                             in_data[229],
                             in_data[587]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [63:0] lut_33_table = 64'b1111111111111111111100111111111100110011001111110000001100000011;
    wire [5:0] lut_33_select = {
                             in_data[396],
                             in_data[100],
                             in_data[318],
                             in_data[207],
                             in_data[204],
                             in_data[39]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [63:0] lut_34_table = 64'b0000111100001111000011110000111100000000000000000000000000000000;
    wire [5:0] lut_34_select = {
                             in_data[292],
                             in_data[413],
                             in_data[76],
                             in_data[681],
                             in_data[756],
                             in_data[113]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [63:0] lut_35_table = 64'b0000000000000011000000000001001000000000001100110000000000110011;
    wire [5:0] lut_35_select = {
                             in_data[190],
                             in_data[14],
                             in_data[209],
                             in_data[418],
                             in_data[92],
                             in_data[590]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [63:0] lut_36_table = 64'b0011001100110000111111111111000000110011001100001111111111110000;
    wire [5:0] lut_36_select = {
                             in_data[642],
                             in_data[652],
                             in_data[370],
                             in_data[367],
                             in_data[571],
                             in_data[727]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [63:0] lut_37_table = 64'b1111100011110000111111101111100011111000111100001111111111111000;
    wire [5:0] lut_37_select = {
                             in_data[22],
                             in_data[611],
                             in_data[482],
                             in_data[399],
                             in_data[478],
                             in_data[134]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [63:0] lut_38_table = 64'b1111111111111111111111101111111011111111111111001011101010101000;
    wire [5:0] lut_38_select = {
                             in_data[119],
                             in_data[429],
                             in_data[445],
                             in_data[491],
                             in_data[570],
                             in_data[487]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [63:0] lut_39_table = 64'b0101011101010101000000000000000001010101010101010000000000000000;
    wire [5:0] lut_39_select = {
                             in_data[666],
                             in_data[215],
                             in_data[114],
                             in_data[404],
                             in_data[336],
                             in_data[328]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [63:0] lut_40_table = 64'b0000000011110000000000001111111000000000111100000010000011111111;
    wire [5:0] lut_40_select = {
                             in_data[364],
                             in_data[173],
                             in_data[326],
                             in_data[603],
                             in_data[5],
                             in_data[25]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [63:0] lut_41_table = 64'b1111101111111010111110111111101111111011111110111111101110111011;
    wire [5:0] lut_41_select = {
                             in_data[210],
                             in_data[452],
                             in_data[473],
                             in_data[462],
                             in_data[345],
                             in_data[174]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [63:0] lut_42_table = 64'b0001000000000000000110011000000011111011111110101111101011111110;
    wire [5:0] lut_42_select = {
                             in_data[238],
                             in_data[548],
                             in_data[598],
                             in_data[380],
                             in_data[635],
                             in_data[500]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [63:0] lut_43_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_43_select = {
                             in_data[271],
                             in_data[138],
                             in_data[454],
                             in_data[307],
                             in_data[66],
                             in_data[91]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [63:0] lut_44_table = 64'b1111111111111111111111111111111111001100110011001100100011001000;
    wire [5:0] lut_44_select = {
                             in_data[578],
                             in_data[672],
                             in_data[551],
                             in_data[640],
                             in_data[95],
                             in_data[137]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [63:0] lut_45_table = 64'b0100010011001100110011001100110001000100110011001100110011001100;
    wire [5:0] lut_45_select = {
                             in_data[373],
                             in_data[451],
                             in_data[694],
                             in_data[671],
                             in_data[299],
                             in_data[460]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [63:0] lut_46_table = 64'b0111011101111111011101110111111100100010001010100010001010100010;
    wire [5:0] lut_46_select = {
                             in_data[509],
                             in_data[170],
                             in_data[750],
                             in_data[744],
                             in_data[261],
                             in_data[540]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [63:0] lut_47_table = 64'b1011000011110000001000000000000011111111111111110000000011111111;
    wire [5:0] lut_47_select = {
                             in_data[297],
                             in_data[70],
                             in_data[633],
                             in_data[288],
                             in_data[474],
                             in_data[83]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [63:0] lut_48_table = 64'b1111000111110001101100001011000011110001111101011011000010110000;
    wire [5:0] lut_48_select = {
                             in_data[751],
                             in_data[184],
                             in_data[117],
                             in_data[303],
                             in_data[245],
                             in_data[651]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [63:0] lut_49_table = 64'b1111111111111111000000000000110011111111111111110000000000000000;
    wire [5:0] lut_49_select = {
                             in_data[421],
                             in_data[375],
                             in_data[163],
                             in_data[664],
                             in_data[534],
                             in_data[56]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [63:0] lut_50_table = 64'b0010001100100011001010110010101000100011001000110010101100101110;
    wire [5:0] lut_50_select = {
                             in_data[306],
                             in_data[604],
                             in_data[277],
                             in_data[268],
                             in_data[458],
                             in_data[627]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [63:0] lut_51_table = 64'b0011001100000001000100110000000100010011000000110001001100010001;
    wire [5:0] lut_51_select = {
                             in_data[589],
                             in_data[213],
                             in_data[305],
                             in_data[547],
                             in_data[566],
                             in_data[740]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [63:0] lut_52_table = 64'b0000111100001111000001010000000010111111001011110000111100000000;
    wire [5:0] lut_52_select = {
                             in_data[165],
                             in_data[572],
                             in_data[126],
                             in_data[638],
                             in_data[31],
                             in_data[423]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [63:0] lut_53_table = 64'b0010101010111111001010101011111100101010101111110010101010111111;
    wire [5:0] lut_53_select = {
                             in_data[7],
                             in_data[667],
                             in_data[300],
                             in_data[564],
                             in_data[466],
                             in_data[192]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [63:0] lut_54_table = 64'b1100110000000000110011001111111111001100000000001100110011111111;
    wire [5:0] lut_54_select = {
                             in_data[23],
                             in_data[313],
                             in_data[543],
                             in_data[6],
                             in_data[537],
                             in_data[29]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [63:0] lut_55_table = 64'b1111111111110000111111111111000011111111111100001111111111110000;
    wire [5:0] lut_55_select = {
                             in_data[255],
                             in_data[15],
                             in_data[637],
                             in_data[527],
                             in_data[18],
                             in_data[467]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [63:0] lut_56_table = 64'b0000111100001111000011110000011101001111000011110000111100001111;
    wire [5:0] lut_56_select = {
                             in_data[729],
                             in_data[217],
                             in_data[106],
                             in_data[461],
                             in_data[759],
                             in_data[757]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [63:0] lut_57_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_57_select = {
                             in_data[726],
                             in_data[146],
                             in_data[595],
                             in_data[242],
                             in_data[617],
                             in_data[650]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [63:0] lut_58_table = 64'b1101110011001100110011000000000011111111111111111100110011001100;
    wire [5:0] lut_58_select = {
                             in_data[395],
                             in_data[158],
                             in_data[350],
                             in_data[533],
                             in_data[463],
                             in_data[778]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [63:0] lut_59_table = 64'b1111111111111111111111111111010101011111010101010101110100000101;
    wire [5:0] lut_59_select = {
                             in_data[655],
                             in_data[704],
                             in_data[746],
                             in_data[187],
                             in_data[777],
                             in_data[372]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [63:0] lut_60_table = 64'b0000000000000000000000000000000011111101111111011111110111111101;
    wire [5:0] lut_60_select = {
                             in_data[220],
                             in_data[703],
                             in_data[646],
                             in_data[665],
                             in_data[705],
                             in_data[291]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [63:0] lut_61_table = 64'b0000001000000010000010100000101000000011000000110000101100001111;
    wire [5:0] lut_61_select = {
                             in_data[630],
                             in_data[290],
                             in_data[96],
                             in_data[247],
                             in_data[136],
                             in_data[544]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [63:0] lut_62_table = 64'b1111111110111010111111101010000011111111111111101111111011101100;
    wire [5:0] lut_62_select = {
                             in_data[680],
                             in_data[497],
                             in_data[539],
                             in_data[360],
                             in_data[409],
                             in_data[455]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [63:0] lut_63_table = 64'b0000000000000000001010100000001000000010000000001011111100101011;
    wire [5:0] lut_63_select = {
                             in_data[609],
                             in_data[686],
                             in_data[102],
                             in_data[175],
                             in_data[384],
                             in_data[591]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [63:0] lut_64_table = 64'b0000000011111111000000001111111100000000111111110000010011111111;
    wire [5:0] lut_64_select = {
                             in_data[45],
                             in_data[448],
                             in_data[457],
                             in_data[89],
                             in_data[619],
                             in_data[382]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [63:0] lut_65_table = 64'b0001000100010001000100010001000100000000000100000001000000010000;
    wire [5:0] lut_65_select = {
                             in_data[185],
                             in_data[200],
                             in_data[21],
                             in_data[499],
                             in_data[162],
                             in_data[249]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [63:0] lut_66_table = 64'b1111111111111111111111001111110011111111111111110111010011110100;
    wire [5:0] lut_66_select = {
                             in_data[13],
                             in_data[573],
                             in_data[323],
                             in_data[122],
                             in_data[568],
                             in_data[765]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [63:0] lut_67_table = 64'b1111111111101110111111111110111011111111110011001111111111001100;
    wire [5:0] lut_67_select = {
                             in_data[214],
                             in_data[391],
                             in_data[410],
                             in_data[28],
                             in_data[149],
                             in_data[695]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [63:0] lut_68_table = 64'b0000111100001111000011110000111100001111000011110000111100001111;
    wire [5:0] lut_68_select = {
                             in_data[586],
                             in_data[782],
                             in_data[109],
                             in_data[516],
                             in_data[260],
                             in_data[67]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [63:0] lut_69_table = 64'b1111111111101110111011101110111011111111111111111111111111101110;
    wire [5:0] lut_69_select = {
                             in_data[65],
                             in_data[709],
                             in_data[441],
                             in_data[309],
                             in_data[284],
                             in_data[206]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [63:0] lut_70_table = 64'b0000000011000000000000001100100011110011111100111111000011110100;
    wire [5:0] lut_70_select = {
                             in_data[658],
                             in_data[582],
                             in_data[581],
                             in_data[327],
                             in_data[439],
                             in_data[280]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [63:0] lut_71_table = 64'b0000000000000000000000000000000000000000000000001111111111111111;
    wire [5:0] lut_71_select = {
                             in_data[623],
                             in_data[684],
                             in_data[530],
                             in_data[764],
                             in_data[732],
                             in_data[758]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [63:0] lut_72_table = 64'b1111111111111100111111111111111111110000111100001111110011110000;
    wire [5:0] lut_72_select = {
                             in_data[536],
                             in_data[262],
                             in_data[507],
                             in_data[324],
                             in_data[484],
                             in_data[86]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [63:0] lut_73_table = 64'b1100000011110000111100001111101111000000111100001111000011111011;
    wire [5:0] lut_73_select = {
                             in_data[82],
                             in_data[339],
                             in_data[234],
                             in_data[105],
                             in_data[246],
                             in_data[776]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [63:0] lut_74_table = 64'b1111111111111111000011110000111111111111111111110000111100001111;
    wire [5:0] lut_74_select = {
                             in_data[583],
                             in_data[254],
                             in_data[335],
                             in_data[317],
                             in_data[169],
                             in_data[702]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [63:0] lut_75_table = 64'b0000000000000000000000000000000000000000000000001111111111111111;
    wire [5:0] lut_75_select = {
                             in_data[201],
                             in_data[440],
                             in_data[256],
                             in_data[775],
                             in_data[59],
                             in_data[0]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [63:0] lut_76_table = 64'b0011000011110000111110111111101100010000010100001111111111111111;
    wire [5:0] lut_76_select = {
                             in_data[610],
                             in_data[401],
                             in_data[69],
                             in_data[358],
                             in_data[639],
                             in_data[406]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [63:0] lut_77_table = 64'b0001000100010001000100010001000100010001000100010001000100010001;
    wire [5:0] lut_77_select = {
                             in_data[196],
                             in_data[281],
                             in_data[62],
                             in_data[673],
                             in_data[325],
                             in_data[739]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [63:0] lut_78_table = 64'b0000000011111111001100110011001100000000111111110011000000110011;
    wire [5:0] lut_78_select = {
                             in_data[225],
                             in_data[653],
                             in_data[579],
                             in_data[369],
                             in_data[405],
                             in_data[12]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [63:0] lut_79_table = 64'b1111011111111111001100001111001111110011001100110111000100110010;
    wire [5:0] lut_79_select = {
                             in_data[212],
                             in_data[593],
                             in_data[492],
                             in_data[257],
                             in_data[720],
                             in_data[180]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [63:0] lut_80_table = 64'b1100111111001111000000000000000011111111111111111111111111111111;
    wire [5:0] lut_80_select = {
                             in_data[520],
                             in_data[741],
                             in_data[670],
                             in_data[381],
                             in_data[773],
                             in_data[387]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [63:0] lut_81_table = 64'b1011001111111011101110111011101100000000000000000010001010100010;
    wire [5:0] lut_81_select = {
                             in_data[183],
                             in_data[710],
                             in_data[49],
                             in_data[390],
                             in_data[108],
                             in_data[584]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [63:0] lut_82_table = 64'b1111110011111101110111011101110111111101111111111101110111011101;
    wire [5:0] lut_82_select = {
                             in_data[222],
                             in_data[514],
                             in_data[11],
                             in_data[453],
                             in_data[693],
                             in_data[265]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [63:0] lut_83_table = 64'b0010111110101111001011111010111100101111111011110010111111101111;
    wire [5:0] lut_83_select = {
                             in_data[647],
                             in_data[733],
                             in_data[178],
                             in_data[379],
                             in_data[293],
                             in_data[714]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [63:0] lut_84_table = 64'b1111111111111010111010101010101011111111111111101111111111101010;
    wire [5:0] lut_84_select = {
                             in_data[721],
                             in_data[592],
                             in_data[311],
                             in_data[442],
                             in_data[93],
                             in_data[518]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [63:0] lut_85_table = 64'b1111111111111111111011110101000111111111111111111010111101000001;
    wire [5:0] lut_85_select = {
                             in_data[4],
                             in_data[386],
                             in_data[181],
                             in_data[523],
                             in_data[17],
                             in_data[270]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [63:0] lut_86_table = 64'b1010101100001111101111111111111100001010000010000000001100000100;
    wire [5:0] lut_86_select = {
                             in_data[398],
                             in_data[272],
                             in_data[486],
                             in_data[535],
                             in_data[68],
                             in_data[351]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [63:0] lut_87_table = 64'b1111111111111111111111111111111111001100110011000100110011001100;
    wire [5:0] lut_87_select = {
                             in_data[713],
                             in_data[392],
                             in_data[577],
                             in_data[575],
                             in_data[371],
                             in_data[37]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [63:0] lut_88_table = 64'b1111111111111111111101111111111111111111000000001111111111110011;
    wire [5:0] lut_88_select = {
                             in_data[343],
                             in_data[243],
                             in_data[607],
                             in_data[538],
                             in_data[754],
                             in_data[283]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [63:0] lut_89_table = 64'b1111111111101111111111111110111011111111111011101111111111101110;
    wire [5:0] lut_89_select = {
                             in_data[161],
                             in_data[251],
                             in_data[626],
                             in_data[3],
                             in_data[687],
                             in_data[624]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [63:0] lut_90_table = 64'b0011001100100000001100000011000000110011111100010011001100110011;
    wire [5:0] lut_90_select = {
                             in_data[266],
                             in_data[237],
                             in_data[239],
                             in_data[295],
                             in_data[377],
                             in_data[674]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [63:0] lut_91_table = 64'b1000101011101111111100001111111111111111111011111111000011111111;
    wire [5:0] lut_91_select = {
                             in_data[301],
                             in_data[231],
                             in_data[211],
                             in_data[596],
                             in_data[475],
                             in_data[417]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [63:0] lut_92_table = 64'b0101000101010001010100010101000101010001010100010101000101010001;
    wire [5:0] lut_92_select = {
                             in_data[1],
                             in_data[61],
                             in_data[139],
                             in_data[508],
                             in_data[41],
                             in_data[342]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [63:0] lut_93_table = 64'b1111111111111111111111111111000011111111111111111111111111110000;
    wire [5:0] lut_93_select = {
                             in_data[55],
                             in_data[770],
                             in_data[218],
                             in_data[471],
                             in_data[226],
                             in_data[110]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [63:0] lut_94_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_94_select = {
                             in_data[422],
                             in_data[341],
                             in_data[781],
                             in_data[143],
                             in_data[616],
                             in_data[554]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [63:0] lut_95_table = 64'b1000000011111111100000001111111100000000111101010000000011110101;
    wire [5:0] lut_95_select = {
                             in_data[679],
                             in_data[731],
                             in_data[289],
                             in_data[154],
                             in_data[449],
                             in_data[456]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [63:0] lut_96_table = 64'b1100111011001100000011000100110011111111111111111010101010101010;
    wire [5:0] lut_96_select = {
                             in_data[552],
                             in_data[347],
                             in_data[32],
                             in_data[150],
                             in_data[632],
                             in_data[321]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [63:0] lut_97_table = 64'b1111111100001111111111111101111110101111000010101010111100001010;
    wire [5:0] lut_97_select = {
                             in_data[416],
                             in_data[279],
                             in_data[378],
                             in_data[495],
                             in_data[762],
                             in_data[657]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [63:0] lut_98_table = 64'b1111111111001100111111111100110011111111110011001111111111001100;
    wire [5:0] lut_98_select = {
                             in_data[362],
                             in_data[614],
                             in_data[524],
                             in_data[314],
                             in_data[219],
                             in_data[71]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [63:0] lut_99_table = 64'b0001000100000001000100010001000000110011000100110011001100110011;
    wire [5:0] lut_99_select = {
                             in_data[388],
                             in_data[763],
                             in_data[51],
                             in_data[755],
                             in_data[156],
                             in_data[75]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [63:0] lut_100_table = 64'b1011101110111011101110111011101110111011101110101011101110111011;
    wire [5:0] lut_100_select = {
                             in_data[74],
                             in_data[385],
                             in_data[562],
                             in_data[697],
                             in_data[357],
                             in_data[567]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [63:0] lut_101_table = 64'b0101111101011111010100000101000001011111010111110101000001010101;
    wire [5:0] lut_101_select = {
                             in_data[46],
                             in_data[103],
                             in_data[698],
                             in_data[135],
                             in_data[8],
                             in_data[621]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [63:0] lut_102_table = 64'b1111000111111011111111111111111100000000000100000001000000010000;
    wire [5:0] lut_102_select = {
                             in_data[541],
                             in_data[668],
                             in_data[641],
                             in_data[479],
                             in_data[769],
                             in_data[682]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [63:0] lut_103_table = 64'b1111111111111111111111111000101011111111111111111111111111101110;
    wire [5:0] lut_103_select = {
                             in_data[675],
                             in_data[618],
                             in_data[120],
                             in_data[588],
                             in_data[363],
                             in_data[447]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [63:0] lut_104_table = 64'b0000000000000000001100000010000000110011001100110011001100110011;
    wire [5:0] lut_104_select = {
                             in_data[235],
                             in_data[52],
                             in_data[411],
                             in_data[558],
                             in_data[287],
                             in_data[140]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [63:0] lut_105_table = 64'b1100110011111111010000001100110011000010111111110000000000000000;
    wire [5:0] lut_105_select = {
                             in_data[496],
                             in_data[244],
                             in_data[715],
                             in_data[553],
                             in_data[127],
                             in_data[194]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [63:0] lut_106_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_106_select = {
                             in_data[515],
                             in_data[737],
                             in_data[636],
                             in_data[87],
                             in_data[227],
                             in_data[688]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [63:0] lut_107_table = 64'b1111101110111010111110111010101011111111111010101111111110101010;
    wire [5:0] lut_107_select = {
                             in_data[50],
                             in_data[768],
                             in_data[188],
                             in_data[498],
                             in_data[772],
                             in_data[240]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [63:0] lut_108_table = 64'b1010101011111111101010101111101110101010111111111010101011111111;
    wire [5:0] lut_108_select = {
                             in_data[569],
                             in_data[716],
                             in_data[349],
                             in_data[476],
                             in_data[532],
                             in_data[202]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [63:0] lut_109_table = 64'b0000000011111111000000000001001100000000001111110000000000000000;
    wire [5:0] lut_109_select = {
                             in_data[722],
                             in_data[691],
                             in_data[556],
                             in_data[36],
                             in_data[72],
                             in_data[115]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [63:0] lut_110_table = 64'b0101010101010100010101010100010101110011001100101111001110110011;
    wire [5:0] lut_110_select = {
                             in_data[469],
                             in_data[734],
                             in_data[133],
                             in_data[597],
                             in_data[438],
                             in_data[273]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [63:0] lut_111_table = 64'b0011011100110011001100110011001100110111001100110011001100110011;
    wire [5:0] lut_111_select = {
                             in_data[308],
                             in_data[124],
                             in_data[259],
                             in_data[315],
                             in_data[430],
                             in_data[253]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [63:0] lut_112_table = 64'b1111111111111111111111110000111111111111111111111111111100000000;
    wire [5:0] lut_112_select = {
                             in_data[278],
                             in_data[660],
                             in_data[118],
                             in_data[121],
                             in_data[615],
                             in_data[90]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [63:0] lut_113_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_113_select = {
                             in_data[493],
                             in_data[85],
                             in_data[81],
                             in_data[282],
                             in_data[157],
                             in_data[80]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [63:0] lut_114_table = 64'b1010111110101011101111111010101110101011101010111011101110101011;
    wire [5:0] lut_114_select = {
                             in_data[224],
                             in_data[78],
                             in_data[248],
                             in_data[230],
                             in_data[654],
                             in_data[153]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [63:0] lut_115_table = 64'b1111111101010101111111110101010111011111010101011111110101010101;
    wire [5:0] lut_115_select = {
                             in_data[198],
                             in_data[752],
                             in_data[258],
                             in_data[10],
                             in_data[761],
                             in_data[376]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [63:0] lut_116_table = 64'b0101010101010101010101010101010101010101010101010100010001000100;
    wire [5:0] lut_116_select = {
                             in_data[112],
                             in_data[27],
                             in_data[30],
                             in_data[559],
                             in_data[685],
                             in_data[275]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [63:0] lut_117_table = 64'b1101110111111111110111011111111111001100010011001100110001001100;
    wire [5:0] lut_117_select = {
                             in_data[546],
                             in_data[760],
                             in_data[550],
                             in_data[723],
                             in_data[594],
                             in_data[557]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [63:0] lut_118_table = 64'b0000010100000101000000000000000011000111111001111110010011100100;
    wire [5:0] lut_118_select = {
                             in_data[612],
                             in_data[542],
                             in_data[780],
                             in_data[274],
                             in_data[177],
                             in_data[182]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [63:0] lut_119_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_119_select = {
                             in_data[645],
                             in_data[519],
                             in_data[412],
                             in_data[700],
                             in_data[285],
                             in_data[450]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [63:0] lut_120_table = 64'b1111111111111111111111011111110011111100111111000001110000001000;
    wire [5:0] lut_120_select = {
                             in_data[425],
                             in_data[241],
                             in_data[743],
                             in_data[205],
                             in_data[383],
                             in_data[9]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [63:0] lut_121_table = 64'b0000101100000011000011110000001100001011000000110000101100000011;
    wire [5:0] lut_121_select = {
                             in_data[644],
                             in_data[57],
                             in_data[38],
                             in_data[464],
                             in_data[676],
                             in_data[366]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [63:0] lut_122_table = 64'b0000000000000000000000000000000011111111010111111111111100010101;
    wire [5:0] lut_122_select = {
                             in_data[233],
                             in_data[643],
                             in_data[264],
                             in_data[503],
                             in_data[599],
                             in_data[748]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [63:0] lut_123_table = 64'b1100111011101111110011101110111111001110111011101100110011101110;
    wire [5:0] lut_123_select = {
                             in_data[712],
                             in_data[669],
                             in_data[329],
                             in_data[199],
                             in_data[468],
                             in_data[708]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [63:0] lut_124_table = 64'b0101010101010101010101010101010101010101010101010101010101010101;
    wire [5:0] lut_124_select = {
                             in_data[319],
                             in_data[312],
                             in_data[145],
                             in_data[683],
                             in_data[477],
                             in_data[354]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [63:0] lut_125_table = 64'b0000000000000000000000000000000011111111111111110000000000000000;
    wire [5:0] lut_125_select = {
                             in_data[555],
                             in_data[344],
                             in_data[656],
                             in_data[747],
                             in_data[563],
                             in_data[250]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [63:0] lut_126_table = 64'b1111010011111111111100001111001111110101111111111111000011110000;
    wire [5:0] lut_126_select = {
                             in_data[47],
                             in_data[735],
                             in_data[661],
                             in_data[711],
                             in_data[24],
                             in_data[197]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [63:0] lut_127_table = 64'b0000000001010101010101010101010100000000000000000101000101010101;
    wire [5:0] lut_127_select = {
                             in_data[263],
                             in_data[159],
                             in_data[613],
                             in_data[48],
                             in_data[505],
                             in_data[625]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [63:0] lut_128_table = 64'b1111101110110010111110111011001011111011101100101111101110110010;
    wire [5:0] lut_128_select = {
                             in_data[34],
                             in_data[443],
                             in_data[525],
                             in_data[631],
                             in_data[407],
                             in_data[356]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [63:0] lut_129_table = 64'b1010101000000000101010100000000011111111000100011111111100010001;
    wire [5:0] lut_129_select = {
                             in_data[189],
                             in_data[88],
                             in_data[348],
                             in_data[730],
                             in_data[517],
                             in_data[346]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [63:0] lut_130_table = 64'b1111111100000000111111111111111111111111000000001111111111001100;
    wire [5:0] lut_130_select = {
                             in_data[257],
                             in_data[433],
                             in_data[659],
                             in_data[16],
                             in_data[144],
                             in_data[766]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [63:0] lut_131_table = 64'b1111111111000100111111111100010011111111111011001111111111101100;
    wire [5:0] lut_131_select = {
                             in_data[417],
                             in_data[172],
                             in_data[689],
                             in_data[641],
                             in_data[410],
                             in_data[743]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [63:0] lut_132_table = 64'b0000000000000000010101010000000000000000000000000101010100000000;
    wire [5:0] lut_132_select = {
                             in_data[32],
                             in_data[103],
                             in_data[521],
                             in_data[194],
                             in_data[419],
                             in_data[693]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [63:0] lut_133_table = 64'b0000000000000000000000000000000000000000000000000000000000110011;
    wire [5:0] lut_133_select = {
                             in_data[509],
                             in_data[129],
                             in_data[122],
                             in_data[649],
                             in_data[127],
                             in_data[82]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [63:0] lut_134_table = 64'b1111111111111111111100111111001111110111111011110100000101000000;
    wire [5:0] lut_134_select = {
                             in_data[552],
                             in_data[191],
                             in_data[101],
                             in_data[602],
                             in_data[578],
                             in_data[549]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [63:0] lut_135_table = 64'b0000111110101111000011110000111100000000001100110000000000100001;
    wire [5:0] lut_135_select = {
                             in_data[655],
                             in_data[604],
                             in_data[398],
                             in_data[405],
                             in_data[107],
                             in_data[454]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [63:0] lut_136_table = 64'b0000000000110011000000000011001100000000010101110000000001111111;
    wire [5:0] lut_136_select = {
                             in_data[275],
                             in_data[138],
                             in_data[494],
                             in_data[363],
                             in_data[382],
                             in_data[514]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [63:0] lut_137_table = 64'b0111011111110111011101111111011101110101111101010000000000000000;
    wire [5:0] lut_137_select = {
                             in_data[350],
                             in_data[440],
                             in_data[446],
                             in_data[577],
                             in_data[355],
                             in_data[407]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [63:0] lut_138_table = 64'b0000000000000000111111111111111100000000000000000000000011111101;
    wire [5:0] lut_138_select = {
                             in_data[348],
                             in_data[159],
                             in_data[330],
                             in_data[478],
                             in_data[187],
                             in_data[222]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [63:0] lut_139_table = 64'b1111111111111100111111111111110000110000001100000011000000110000;
    wire [5:0] lut_139_select = {
                             in_data[459],
                             in_data[169],
                             in_data[105],
                             in_data[346],
                             in_data[682],
                             in_data[111]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [63:0] lut_140_table = 64'b0000000000000000000000000000000000000100000000001101110101010101;
    wire [5:0] lut_140_select = {
                             in_data[125],
                             in_data[227],
                             in_data[43],
                             in_data[112],
                             in_data[722],
                             in_data[277]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [63:0] lut_141_table = 64'b0000000000000000000000000000000000000000000000001111100011111111;
    wire [5:0] lut_141_select = {
                             in_data[607],
                             in_data[550],
                             in_data[768],
                             in_data[268],
                             in_data[49],
                             in_data[751]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [63:0] lut_142_table = 64'b1111000011110000111100001111000011110010111100101111001011110010;
    wire [5:0] lut_142_select = {
                             in_data[210],
                             in_data[67],
                             in_data[51],
                             in_data[519],
                             in_data[628],
                             in_data[412]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [63:0] lut_143_table = 64'b0000100000001000000010100000101010001111100011111000111110001111;
    wire [5:0] lut_143_select = {
                             in_data[713],
                             in_data[143],
                             in_data[195],
                             in_data[538],
                             in_data[192],
                             in_data[276]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [63:0] lut_144_table = 64'b1101110111001101110111111100110111001111110011011100111111001101;
    wire [5:0] lut_144_select = {
                             in_data[301],
                             in_data[531],
                             in_data[364],
                             in_data[124],
                             in_data[706],
                             in_data[623]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [63:0] lut_145_table = 64'b0000001000000000001100110011001100111111001111111111111110111111;
    wire [5:0] lut_145_select = {
                             in_data[597],
                             in_data[598],
                             in_data[36],
                             in_data[564],
                             in_data[240],
                             in_data[366]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [63:0] lut_146_table = 64'b1011111100100010111111111011111100101010000000001011111100000010;
    wire [5:0] lut_146_select = {
                             in_data[500],
                             in_data[736],
                             in_data[344],
                             in_data[85],
                             in_data[735],
                             in_data[118]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [63:0] lut_147_table = 64'b0000000000000000001000000000000000000000000000000011001100110011;
    wire [5:0] lut_147_select = {
                             in_data[283],
                             in_data[90],
                             in_data[116],
                             in_data[753],
                             in_data[762],
                             in_data[698]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [63:0] lut_148_table = 64'b1111000011110000111111101111110011110000111100001111000011110000;
    wire [5:0] lut_148_select = {
                             in_data[428],
                             in_data[207],
                             in_data[445],
                             in_data[455],
                             in_data[477],
                             in_data[223]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [63:0] lut_149_table = 64'b0101010111111111011101011111011101010101011101010101010001110101;
    wire [5:0] lut_149_select = {
                             in_data[77],
                             in_data[763],
                             in_data[400],
                             in_data[525],
                             in_data[236],
                             in_data[465]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [63:0] lut_150_table = 64'b0011111100111111001111110000001100111111000100110011001100000000;
    wire [5:0] lut_150_select = {
                             in_data[453],
                             in_data[183],
                             in_data[594],
                             in_data[320],
                             in_data[100],
                             in_data[367]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [63:0] lut_151_table = 64'b1111010111110101111101011111010111110101111101011111010011110101;
    wire [5:0] lut_151_select = {
                             in_data[390],
                             in_data[420],
                             in_data[12],
                             in_data[273],
                             in_data[337],
                             in_data[186]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [63:0] lut_152_table = 64'b0011001000100000101100110010001010110011001100101011101100110011;
    wire [5:0] lut_152_select = {
                             in_data[738],
                             in_data[451],
                             in_data[640],
                             in_data[74],
                             in_data[220],
                             in_data[136]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [63:0] lut_153_table = 64'b0011000011110010001100000000000000110010111111111111001111110111;
    wire [5:0] lut_153_select = {
                             in_data[461],
                             in_data[151],
                             in_data[485],
                             in_data[165],
                             in_data[721],
                             in_data[254]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [63:0] lut_154_table = 64'b0001000000000000000100000000000000010101000000000101010100000100;
    wire [5:0] lut_154_select = {
                             in_data[584],
                             in_data[260],
                             in_data[324],
                             in_data[299],
                             in_data[234],
                             in_data[583]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [63:0] lut_155_table = 64'b0000000010100000000000001010000010101010111110101010101011111010;
    wire [5:0] lut_155_select = {
                             in_data[650],
                             in_data[18],
                             in_data[131],
                             in_data[161],
                             in_data[671],
                             in_data[319]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [63:0] lut_156_table = 64'b1000100011111111100000001111111100000000000000000000000000010000;
    wire [5:0] lut_156_select = {
                             in_data[486],
                             in_data[25],
                             in_data[188],
                             in_data[84],
                             in_data[632],
                             in_data[568]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [63:0] lut_157_table = 64'b1111111111111111000001011111111100000000000000000000000000000000;
    wire [5:0] lut_157_select = {
                             in_data[378],
                             in_data[269],
                             in_data[388],
                             in_data[360],
                             in_data[696],
                             in_data[467]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [63:0] lut_158_table = 64'b0100000000000000000000000000000000001111110011110000111100001111;
    wire [5:0] lut_158_select = {
                             in_data[300],
                             in_data[8],
                             in_data[776],
                             in_data[289],
                             in_data[387],
                             in_data[562]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [63:0] lut_159_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_159_select = {
                             in_data[152],
                             in_data[23],
                             in_data[353],
                             in_data[755],
                             in_data[517],
                             in_data[57]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [63:0] lut_160_table = 64'b0000000000000000101010101010000010101010101010101111101011111110;
    wire [5:0] lut_160_select = {
                             in_data[690],
                             in_data[371],
                             in_data[427],
                             in_data[647],
                             in_data[560],
                             in_data[380]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [63:0] lut_161_table = 64'b1110111011101110111111111111111111101110111011101111111011111111;
    wire [5:0] lut_161_select = {
                             in_data[757],
                             in_data[600],
                             in_data[312],
                             in_data[396],
                             in_data[190],
                             in_data[694]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [63:0] lut_162_table = 64'b0000000011001100000110011100110000000000110011000001100111001100;
    wire [5:0] lut_162_select = {
                             in_data[644],
                             in_data[677],
                             in_data[544],
                             in_data[339],
                             in_data[401],
                             in_data[354]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [63:0] lut_163_table = 64'b1111000010110000111110101111101011111111010100001111111111110101;
    wire [5:0] lut_163_select = {
                             in_data[466],
                             in_data[711],
                             in_data[158],
                             in_data[150],
                             in_data[45],
                             in_data[553]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [63:0] lut_164_table = 64'b0000111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_164_select = {
                             in_data[94],
                             in_data[515],
                             in_data[452],
                             in_data[267],
                             in_data[619],
                             in_data[29]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [63:0] lut_165_table = 64'b0000000000000000000011001111110000001111000000000000111111111100;
    wire [5:0] lut_165_select = {
                             in_data[237],
                             in_data[416],
                             in_data[574],
                             in_data[239],
                             in_data[590],
                             in_data[221]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [63:0] lut_166_table = 64'b0101010101010101010001000100010001010101010101010000010000000100;
    wire [5:0] lut_166_select = {
                             in_data[64],
                             in_data[464],
                             in_data[617],
                             in_data[147],
                             in_data[432],
                             in_data[679]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [63:0] lut_167_table = 64'b0000000000000101000000001111010100000000000001010000000011110101;
    wire [5:0] lut_167_select = {
                             in_data[724],
                             in_data[572],
                             in_data[153],
                             in_data[285],
                             in_data[206],
                             in_data[471]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [63:0] lut_168_table = 64'b1110111111101111111011111110111111101111111011111110111111101111;
    wire [5:0] lut_168_select = {
                             in_data[727],
                             in_data[114],
                             in_data[702],
                             in_data[386],
                             in_data[712],
                             in_data[744]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [63:0] lut_169_table = 64'b1111111111111111111011101110111011111111111111111110111011101110;
    wire [5:0] lut_169_select = {
                             in_data[27],
                             in_data[566],
                             in_data[309],
                             in_data[139],
                             in_data[506],
                             in_data[444]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [63:0] lut_170_table = 64'b0001011100010101001111110001010111011101000101011101110100000101;
    wire [5:0] lut_170_select = {
                             in_data[493],
                             in_data[771],
                             in_data[304],
                             in_data[536],
                             in_data[245],
                             in_data[545]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [63:0] lut_171_table = 64'b0000101000001111000010100000111100000010000011110000101000001111;
    wire [5:0] lut_171_select = {
                             in_data[764],
                             in_data[55],
                             in_data[695],
                             in_data[662],
                             in_data[646],
                             in_data[342]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [63:0] lut_172_table = 64'b1000100000000000000000001111111100000000000000000000000011111111;
    wire [5:0] lut_172_select = {
                             in_data[576],
                             in_data[97],
                             in_data[208],
                             in_data[672],
                             in_data[608],
                             in_data[133]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [63:0] lut_173_table = 64'b1111111111111111111111111111111111110000111100001111000011110000;
    wire [5:0] lut_173_select = {
                             in_data[431],
                             in_data[88],
                             in_data[703],
                             in_data[93],
                             in_data[612],
                             in_data[219]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [63:0] lut_174_table = 64'b1111101011111011111111111111111100000000000000000001000000010000;
    wire [5:0] lut_174_select = {
                             in_data[434],
                             in_data[154],
                             in_data[137],
                             in_data[331],
                             in_data[306],
                             in_data[481]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [63:0] lut_175_table = 64'b1100110011001100110011111100111111001100110011001100111011001100;
    wire [5:0] lut_175_select = {
                             in_data[228],
                             in_data[415],
                             in_data[395],
                             in_data[516],
                             in_data[266],
                             in_data[653]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [63:0] lut_176_table = 64'b1111111111110111110101110101010111111111011101010101010101010101;
    wire [5:0] lut_176_select = {
                             in_data[79],
                             in_data[134],
                             in_data[535],
                             in_data[7],
                             in_data[59],
                             in_data[687]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [63:0] lut_177_table = 64'b1110111111111111110011111110111111001111100011111100111010001110;
    wire [5:0] lut_177_select = {
                             in_data[274],
                             in_data[534],
                             in_data[651],
                             in_data[294],
                             in_data[205],
                             in_data[120]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [63:0] lut_178_table = 64'b0000000000000000000000000000000000010001000100000000101000001010;
    wire [5:0] lut_178_select = {
                             in_data[593],
                             in_data[209],
                             in_data[50],
                             in_data[264],
                             in_data[175],
                             in_data[462]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [63:0] lut_179_table = 64'b0100010101000100010001000100010001000100010011000100010001000101;
    wire [5:0] lut_179_select = {
                             in_data[372],
                             in_data[335],
                             in_data[501],
                             in_data[758],
                             in_data[626],
                             in_data[463]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [63:0] lut_180_table = 64'b0000000000000000000000001011111100000000000000000000000011111111;
    wire [5:0] lut_180_select = {
                             in_data[760],
                             in_data[326],
                             in_data[162],
                             in_data[216],
                             in_data[767],
                             in_data[393]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [63:0] lut_181_table = 64'b0011001100110011001100110011000100110011001100110011001100110011;
    wire [5:0] lut_181_select = {
                             in_data[19],
                             in_data[730],
                             in_data[213],
                             in_data[476],
                             in_data[606],
                             in_data[76]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [63:0] lut_182_table = 64'b1110110000000000111111111111111111001100000000001111111011111111;
    wire [5:0] lut_182_select = {
                             in_data[773],
                             in_data[316],
                             in_data[343],
                             in_data[614],
                             in_data[265],
                             in_data[561]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [63:0] lut_183_table = 64'b1100110011001100110011011100110100000000000000000000000000000001;
    wire [5:0] lut_183_select = {
                             in_data[297],
                             in_data[551],
                             in_data[253],
                             in_data[480],
                             in_data[375],
                             in_data[149]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [63:0] lut_184_table = 64'b1111111110100101101011110000000011111111000001011010111100000101;
    wire [5:0] lut_184_select = {
                             in_data[504],
                             in_data[648],
                             in_data[484],
                             in_data[376],
                             in_data[505],
                             in_data[457]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [63:0] lut_185_table = 64'b1100110011001100111111111111111111001100110011001100110011001100;
    wire [5:0] lut_185_select = {
                             in_data[66],
                             in_data[527],
                             in_data[352],
                             in_data[700],
                             in_data[414],
                             in_data[587]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [63:0] lut_186_table = 64'b0000000000000000000000000101010100000000000000000000000001010101;
    wire [5:0] lut_186_select = {
                             in_data[40],
                             in_data[745],
                             in_data[585],
                             in_data[307],
                             in_data[141],
                             in_data[438]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [63:0] lut_187_table = 64'b1111111111111111111111111111000011111111111111111111111111111001;
    wire [5:0] lut_187_select = {
                             in_data[252],
                             in_data[75],
                             in_data[557],
                             in_data[479],
                             in_data[196],
                             in_data[52]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [63:0] lut_188_table = 64'b1000000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_188_select = {
                             in_data[166],
                             in_data[176],
                             in_data[765],
                             in_data[513],
                             in_data[613],
                             in_data[365]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [63:0] lut_189_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_189_select = {
                             in_data[171],
                             in_data[261],
                             in_data[63],
                             in_data[547],
                             in_data[756],
                             in_data[413]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [63:0] lut_190_table = 64'b0101010101010101010101010101010101000101000000000101010101010101;
    wire [5:0] lut_190_select = {
                             in_data[246],
                             in_data[656],
                             in_data[9],
                             in_data[769],
                             in_data[759],
                             in_data[439]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [63:0] lut_191_table = 64'b0000000000000000000000000000000000000000011111110000000001111111;
    wire [5:0] lut_191_select = {
                             in_data[119],
                             in_data[35],
                             in_data[290],
                             in_data[115],
                             in_data[197],
                             in_data[422]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [63:0] lut_192_table = 64'b1111111101010100111111110101010011111111010001011111111101010101;
    wire [5:0] lut_192_select = {
                             in_data[603],
                             in_data[383],
                             in_data[146],
                             in_data[615],
                             in_data[775],
                             in_data[660]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [63:0] lut_193_table = 64'b0000000001010101000000000101010100000000010101010000000001010101;
    wire [5:0] lut_193_select = {
                             in_data[24],
                             in_data[643],
                             in_data[262],
                             in_data[750],
                             in_data[89],
                             in_data[739]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [63:0] lut_194_table = 64'b1111111111111111111111111111111111111111111111111111000011111000;
    wire [5:0] lut_194_select = {
                             in_data[621],
                             in_data[126],
                             in_data[323],
                             in_data[567],
                             in_data[148],
                             in_data[697]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [63:0] lut_195_table = 64'b0000000001010101010001010101010100000000010101010000010001010101;
    wire [5:0] lut_195_select = {
                             in_data[22],
                             in_data[53],
                             in_data[540],
                             in_data[81],
                             in_data[20],
                             in_data[683]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [63:0] lut_196_table = 64'b1111111100110011111111110000000011111111001100111100110000000000;
    wire [5:0] lut_196_select = {
                             in_data[473],
                             in_data[322],
                             in_data[314],
                             in_data[46],
                             in_data[634],
                             in_data[3]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [63:0] lut_197_table = 64'b1111110111001100111111111111110111110101110100001111110111110000;
    wire [5:0] lut_197_select = {
                             in_data[498],
                             in_data[332],
                             in_data[620],
                             in_data[179],
                             in_data[347],
                             in_data[385]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [63:0] lut_198_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_198_select = {
                             in_data[145],
                             in_data[255],
                             in_data[408],
                             in_data[113],
                             in_data[315],
                             in_data[539]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [63:0] lut_199_table = 64'b0000000000000000000011110000000001001111010001001111111100001101;
    wire [5:0] lut_199_select = {
                             in_data[70],
                             in_data[573],
                             in_data[303],
                             in_data[678],
                             in_data[204],
                             in_data[328]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [63:0] lut_200_table = 64'b0001001100110011001100110011001100000011000100110000001100010011;
    wire [5:0] lut_200_select = {
                             in_data[44],
                             in_data[726],
                             in_data[167],
                             in_data[708],
                             in_data[605],
                             in_data[394]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [63:0] lut_201_table = 64'b1100000011111100110011001111110011000000111111001100110011111100;
    wire [5:0] lut_201_select = {
                             in_data[110],
                             in_data[281],
                             in_data[748],
                             in_data[42],
                             in_data[201],
                             in_data[674]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [63:0] lut_202_table = 64'b0000101000100010001010100010101100001110001011110010111000101111;
    wire [5:0] lut_202_select = {
                             in_data[135],
                             in_data[482],
                             in_data[123],
                             in_data[520],
                             in_data[524],
                             in_data[259]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [63:0] lut_203_table = 64'b1111000111111111111100001111111101010000111100000101000011110000;
    wire [5:0] lut_203_select = {
                             in_data[178],
                             in_data[533],
                             in_data[510],
                             in_data[241],
                             in_data[443],
                             in_data[218]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [63:0] lut_204_table = 64'b0011001000110010001000100010001000110010001100100011001000110010;
    wire [5:0] lut_204_select = {
                             in_data[117],
                             in_data[98],
                             in_data[1],
                             in_data[460],
                             in_data[507],
                             in_data[349]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [63:0] lut_205_table = 64'b0000000000000000001100110011001100000000000000000011001100110011;
    wire [5:0] lut_205_select = {
                             in_data[142],
                             in_data[302],
                             in_data[174],
                             in_data[667],
                             in_data[272],
                             in_data[638]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [63:0] lut_206_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_206_select = {
                             in_data[226],
                             in_data[670],
                             in_data[327],
                             in_data[95],
                             in_data[686],
                             in_data[106]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [63:0] lut_207_table = 64'b1111000011111110100000001011111111100000111111010000000011011111;
    wire [5:0] lut_207_select = {
                             in_data[778],
                             in_data[321],
                             in_data[406],
                             in_data[488],
                             in_data[503],
                             in_data[78]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [63:0] lut_208_table = 64'b1010101010101000111111111111101010101010101010101111111111111111;
    wire [5:0] lut_208_select = {
                             in_data[173],
                             in_data[496],
                             in_data[546],
                             in_data[305],
                             in_data[10],
                             in_data[716]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [63:0] lut_209_table = 64'b1110111111111111111011111110111111001100111011101000111010101110;
    wire [5:0] lut_209_select = {
                             in_data[442],
                             in_data[637],
                             in_data[747],
                             in_data[68],
                             in_data[359],
                             in_data[155]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [63:0] lut_210_table = 64'b0000000100000101000000110000001100000001000001010000001100000011;
    wire [5:0] lut_210_select = {
                             in_data[13],
                             in_data[652],
                             in_data[15],
                             in_data[497],
                             in_data[73],
                             in_data[625]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [63:0] lut_211_table = 64'b1111111111111111111111101111111111101100111011001110110011101100;
    wire [5:0] lut_211_select = {
                             in_data[373],
                             in_data[170],
                             in_data[624],
                             in_data[468],
                             in_data[329],
                             in_data[357]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [63:0] lut_212_table = 64'b0000000001111111000000000011111100000000000111110000000000001111;
    wire [5:0] lut_212_select = {
                             in_data[421],
                             in_data[224],
                             in_data[458],
                             in_data[230],
                             in_data[308],
                             in_data[58]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [63:0] lut_213_table = 64'b1111111111111111111111111100110011111111111111111110110111001100;
    wire [5:0] lut_213_select = {
                             in_data[669],
                             in_data[436],
                             in_data[774],
                             in_data[30],
                             in_data[668],
                             in_data[26]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [63:0] lut_214_table = 64'b0000000000000111000001010101010100000000000001010000010101000101;
    wire [5:0] lut_214_select = {
                             in_data[725],
                             in_data[180],
                             in_data[592],
                             in_data[489],
                             in_data[65],
                             in_data[635]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [63:0] lut_215_table = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    wire [5:0] lut_215_select = {
                             in_data[714],
                             in_data[229],
                             in_data[636],
                             in_data[718],
                             in_data[588],
                             in_data[589]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [63:0] lut_216_table = 64'b0100000011000000110100001101000001000000010000000101000011010000;
    wire [5:0] lut_216_select = {
                             in_data[244],
                             in_data[313],
                             in_data[336],
                             in_data[379],
                             in_data[325],
                             in_data[742]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [63:0] lut_217_table = 64'b1111111111111111110111111111111111011101110011010000000010000000;
    wire [5:0] lut_217_select = {
                             in_data[580],
                             in_data[399],
                             in_data[542],
                             in_data[475],
                             in_data[575],
                             in_data[163]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [63:0] lut_218_table = 64'b0010001100100011001000110010001100000010001000110000001100100011;
    wire [5:0] lut_218_select = {
                             in_data[618],
                             in_data[160],
                             in_data[80],
                             in_data[263],
                             in_data[341],
                             in_data[491]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [63:0] lut_219_table = 64'b1111111111111111111111111111111111111111000000000000000000000000;
    wire [5:0] lut_219_select = {
                             in_data[570],
                             in_data[291],
                             in_data[554],
                             in_data[38],
                             in_data[779],
                             in_data[0]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [63:0] lut_220_table = 64'b0000000000000000000000000001000100000000001100110000000000110011;
    wire [5:0] lut_220_select = {
                             in_data[402],
                             in_data[437],
                             in_data[121],
                             in_data[391],
                             in_data[555],
                             in_data[599]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [63:0] lut_221_table = 64'b0000000001111111000000000101111100001010111111110000101011111111;
    wire [5:0] lut_221_select = {
                             in_data[610],
                             in_data[729],
                             in_data[404],
                             in_data[581],
                             in_data[21],
                             in_data[203]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [63:0] lut_222_table = 64'b0000111000001111000011110000111100001110000011110000111100001111;
    wire [5:0] lut_222_select = {
                             in_data[2],
                             in_data[782],
                             in_data[537],
                             in_data[374],
                             in_data[772],
                             in_data[17]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [63:0] lut_223_table = 64'b1101111111011111110111111111111101001101010011010100110101001101;
    wire [5:0] lut_223_select = {
                             in_data[663],
                             in_data[397],
                             in_data[701],
                             in_data[425],
                             in_data[368],
                             in_data[430]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [63:0] lut_224_table = 64'b1111111111111111111101010101111100000000010101010000000000000101;
    wire [5:0] lut_224_select = {
                             in_data[270],
                             in_data[746],
                             in_data[495],
                             in_data[661],
                             in_data[699],
                             in_data[411]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [63:0] lut_225_table = 64'b0000000000000000000001000000000000000000000000000101110101010101;
    wire [5:0] lut_225_select = {
                             in_data[715],
                             in_data[633],
                             in_data[609],
                             in_data[389],
                             in_data[733],
                             in_data[657]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [63:0] lut_226_table = 64'b0011001011111111001100000011000000111111001111110011000000111100;
    wire [5:0] lut_226_select = {
                             in_data[492],
                             in_data[69],
                             in_data[601],
                             in_data[571],
                             in_data[189],
                             in_data[731]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [63:0] lut_227_table = 64'b0000000000000000111111110000000000000000000000001111111111101110;
    wire [5:0] lut_227_select = {
                             in_data[248],
                             in_data[472],
                             in_data[470],
                             in_data[777],
                             in_data[616],
                             in_data[704]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [63:0] lut_228_table = 64'b1100111100000100110011110000010011001100110011001100110011001100;
    wire [5:0] lut_228_select = {
                             in_data[522],
                             in_data[447],
                             in_data[217],
                             in_data[286],
                             in_data[185],
                             in_data[737]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [63:0] lut_229_table = 64'b1111111111111111111010001111111011111111111111111010100011101000;
    wire [5:0] lut_229_select = {
                             in_data[734],
                             in_data[345],
                             in_data[5],
                             in_data[242],
                             in_data[665],
                             in_data[666]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [63:0] lut_230_table = 64'b0101111111111110010111111111111110101010101010100111111110101010;
    wire [5:0] lut_230_select = {
                             in_data[543],
                             in_data[6],
                             in_data[156],
                             in_data[298],
                             in_data[56],
                             in_data[177]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [63:0] lut_231_table = 64'b1111111111111111111111111111111011111111111111111111111111111010;
    wire [5:0] lut_231_select = {
                             in_data[250],
                             in_data[310],
                             in_data[99],
                             in_data[681],
                             in_data[559],
                             in_data[157]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [63:0] lut_232_table = 64'b1111111100110011111111110011001100110011000000000011001100000000;
    wire [5:0] lut_232_select = {
                             in_data[381],
                             in_data[392],
                             in_data[361],
                             in_data[34],
                             in_data[654],
                             in_data[675]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [63:0] lut_233_table = 64'b1010000011101111101000001110111110100000111011111010000011101111;
    wire [5:0] lut_233_select = {
                             in_data[450],
                             in_data[62],
                             in_data[296],
                             in_data[258],
                             in_data[369],
                             in_data[370]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [63:0] lut_234_table = 64'b0000000000000000111111111111111100000000000000001111111101110111;
    wire [5:0] lut_234_select = {
                             in_data[639],
                             in_data[128],
                             in_data[271],
                             in_data[783],
                             in_data[732],
                             in_data[251]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [63:0] lut_235_table = 64'b1111001111010000111101111111110110010000111111001111000111111101;
    wire [5:0] lut_235_select = {
                             in_data[490],
                             in_data[92],
                             in_data[293],
                             in_data[719],
                             in_data[232],
                             in_data[351]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [63:0] lut_236_table = 64'b0000110000001100000011100000111000001100000011100000111000001110;
    wire [5:0] lut_236_select = {
                             in_data[47],
                             in_data[426],
                             in_data[362],
                             in_data[132],
                             in_data[658],
                             in_data[284]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [63:0] lut_237_table = 64'b1101110111011101110100011101000111011101110110011001000100010001;
    wire [5:0] lut_237_select = {
                             in_data[508],
                             in_data[181],
                             in_data[645],
                             in_data[595],
                             in_data[403],
                             in_data[429]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [63:0] lut_238_table = 64'b0011111100000011001111110000001100100011000000000011001100000011;
    wire [5:0] lut_238_select = {
                             in_data[680],
                             in_data[423],
                             in_data[740],
                             in_data[596],
                             in_data[622],
                             in_data[33]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [63:0] lut_239_table = 64'b1111111111111111111111111111111111111000111111001111100011111000;
    wire [5:0] lut_239_select = {
                             in_data[691],
                             in_data[14],
                             in_data[676],
                             in_data[231],
                             in_data[424],
                             in_data[249]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [63:0] lut_240_table = 64'b1110101110001011101000000000000000000011000011110000000000000011;
    wire [5:0] lut_240_select = {
                             in_data[526],
                             in_data[685],
                             in_data[579],
                             in_data[377],
                             in_data[499],
                             in_data[96]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [63:0] lut_241_table = 64'b0001100100001111111111111111111100001111000011110000111100001111;
    wire [5:0] lut_241_select = {
                             in_data[130],
                             in_data[435],
                             in_data[512],
                             in_data[238],
                             in_data[61],
                             in_data[532]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [63:0] lut_242_table = 64'b0000000000000000000000000000000011111111111111011111111111111101;
    wire [5:0] lut_242_select = {
                             in_data[182],
                             in_data[198],
                             in_data[629],
                             in_data[41],
                             in_data[48],
                             in_data[754]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [63:0] lut_243_table = 64'b0000000000000000000000000000000000000000000000001100010011001100;
    wire [5:0] lut_243_select = {
                             in_data[556],
                             in_data[282],
                             in_data[54],
                             in_data[109],
                             in_data[211],
                             in_data[529]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [63:0] lut_244_table = 64'b1111111011111111111111011111110111101000111111101101110111111101;
    wire [5:0] lut_244_select = {
                             in_data[528],
                             in_data[215],
                             in_data[591],
                             in_data[288],
                             in_data[611],
                             in_data[630]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [63:0] lut_245_table = 64'b0000000000000000000000000000000001010101010101010101010101010101;
    wire [5:0] lut_245_select = {
                             in_data[317],
                             in_data[781],
                             in_data[83],
                             in_data[723],
                             in_data[563],
                             in_data[692]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [63:0] lut_246_table = 64'b1111111100000000101111111010101011111111000000001111111111111010;
    wire [5:0] lut_246_select = {
                             in_data[409],
                             in_data[688],
                             in_data[684],
                             in_data[334],
                             in_data[87],
                             in_data[243]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [63:0] lut_247_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_247_select = {
                             in_data[247],
                             in_data[474],
                             in_data[642],
                             in_data[340],
                             in_data[212],
                             in_data[780]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [63:0] lut_248_table = 64'b1111111101110101111101110101000011111111111111110101000000000000;
    wire [5:0] lut_248_select = {
                             in_data[523],
                             in_data[318],
                             in_data[311],
                             in_data[338],
                             in_data[86],
                             in_data[91]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [63:0] lut_249_table = 64'b1111111111111111111111111111101011111111111111111111111111111010;
    wire [5:0] lut_249_select = {
                             in_data[225],
                             in_data[418],
                             in_data[720],
                             in_data[358],
                             in_data[279],
                             in_data[72]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [63:0] lut_250_table = 64'b1010101010111011101010101010101010111011101111111011101110111011;
    wire [5:0] lut_250_select = {
                             in_data[627],
                             in_data[502],
                             in_data[749],
                             in_data[60],
                             in_data[356],
                             in_data[256]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [63:0] lut_251_table = 64'b0000000000000000000000000000000000010000000100000000010100000101;
    wire [5:0] lut_251_select = {
                             in_data[202],
                             in_data[384],
                             in_data[11],
                             in_data[469],
                             in_data[586],
                             in_data[770]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [63:0] lut_252_table = 64'b1111111100001111111111110000111111111111000011111111111100001111;
    wire [5:0] lut_252_select = {
                             in_data[448],
                             in_data[37],
                             in_data[287],
                             in_data[631],
                             in_data[199],
                             in_data[280]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [63:0] lut_253_table = 64'b0101010100000000000101010000000001010101000000000101010100000000;
    wire [5:0] lut_253_select = {
                             in_data[200],
                             in_data[728],
                             in_data[518],
                             in_data[193],
                             in_data[333],
                             in_data[292]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [63:0] lut_254_table = 64'b1111111111110101111111111111011111110000111100001111010111110000;
    wire [5:0] lut_254_select = {
                             in_data[295],
                             in_data[108],
                             in_data[709],
                             in_data[565],
                             in_data[752],
                             in_data[541]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [63:0] lut_255_table = 64'b1010111100000010111111110010001110101111000000101111111100100011;
    wire [5:0] lut_255_select = {
                             in_data[449],
                             in_data[483],
                             in_data[441],
                             in_data[511],
                             in_data[184],
                             in_data[664]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [63:0] lut_256_table = 64'b1111111111111111111111111111110011111111111111111111111111111100;
    wire [5:0] lut_256_select = {
                             in_data[4],
                             in_data[104],
                             in_data[707],
                             in_data[530],
                             in_data[102],
                             in_data[761]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [63:0] lut_257_table = 64'b1111111110101010111111111010101011111111111110101111111111101010;
    wire [5:0] lut_257_select = {
                             in_data[71],
                             in_data[741],
                             in_data[233],
                             in_data[582],
                             in_data[28],
                             in_data[456]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [63:0] lut_258_table = 64'b1111011100110011111101110011001111110011001100111111111100110011;
    wire [5:0] lut_258_select = {
                             in_data[140],
                             in_data[673],
                             in_data[558],
                             in_data[39],
                             in_data[214],
                             in_data[31]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [63:0] lut_259_table = 64'b0010001011101110000000001010111000100010101010100010000010101010;
    wire [5:0] lut_259_select = {
                             in_data[235],
                             in_data[164],
                             in_data[710],
                             in_data[278],
                             in_data[717],
                             in_data[548]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [63:0] lut_260_table = 64'b0000110011001111000011000000110000001100000011110000110000001100;
    wire [5:0] lut_260_select = {
                             in_data[43],
                             in_data[103],
                             in_data[487],
                             in_data[705],
                             in_data[569],
                             in_data[168]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [63:0] lut_261_table = 64'b1111111111111111111111111111111011000000111010001000000011101000;
    wire [5:0] lut_261_select = {
                             in_data[295],
                             in_data[668],
                             in_data[220],
                             in_data[529],
                             in_data[267],
                             in_data[70]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [63:0] lut_262_table = 64'b0111011100110000001100110010000001110111001100000111001100100000;
    wire [5:0] lut_262_select = {
                             in_data[16],
                             in_data[161],
                             in_data[235],
                             in_data[602],
                             in_data[303],
                             in_data[541]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [63:0] lut_263_table = 64'b1111111100111011111111110011001111111111001100111111111100110011;
    wire [5:0] lut_263_select = {
                             in_data[479],
                             in_data[87],
                             in_data[150],
                             in_data[727],
                             in_data[408],
                             in_data[737]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [63:0] lut_264_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_264_select = {
                             in_data[297],
                             in_data[642],
                             in_data[556],
                             in_data[459],
                             in_data[441],
                             in_data[421]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [63:0] lut_265_table = 64'b0000000000000000000000001111000000000000000000000000000000110000;
    wire [5:0] lut_265_select = {
                             in_data[694],
                             in_data[107],
                             in_data[473],
                             in_data[600],
                             in_data[733],
                             in_data[57]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [63:0] lut_266_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_266_select = {
                             in_data[690],
                             in_data[632],
                             in_data[587],
                             in_data[423],
                             in_data[469],
                             in_data[588]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [63:0] lut_267_table = 64'b0000000011111111000000001010101000001111111111110000000011111111;
    wire [5:0] lut_267_select = {
                             in_data[164],
                             in_data[597],
                             in_data[346],
                             in_data[79],
                             in_data[59],
                             in_data[240]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [63:0] lut_268_table = 64'b0000000000000100000000000000010011001101110011111100111111001111;
    wire [5:0] lut_268_select = {
                             in_data[717],
                             in_data[503],
                             in_data[641],
                             in_data[686],
                             in_data[679],
                             in_data[306]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [63:0] lut_269_table = 64'b0010000000000000001000000000000011110010111100001111001111110010;
    wire [5:0] lut_269_select = {
                             in_data[552],
                             in_data[144],
                             in_data[222],
                             in_data[596],
                             in_data[121],
                             in_data[291]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [63:0] lut_270_table = 64'b0000000000000000000000000000010000000000100011001000100011111111;
    wire [5:0] lut_270_select = {
                             in_data[286],
                             in_data[230],
                             in_data[464],
                             in_data[615],
                             in_data[661],
                             in_data[8]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [63:0] lut_271_table = 64'b0000010100000101000001010000010100000101000001010000010100000101;
    wire [5:0] lut_271_select = {
                             in_data[532],
                             in_data[45],
                             in_data[47],
                             in_data[652],
                             in_data[765],
                             in_data[125]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [63:0] lut_272_table = 64'b1111111111111111010101111111111101000101000000000000000100000000;
    wire [5:0] lut_272_select = {
                             in_data[659],
                             in_data[380],
                             in_data[126],
                             in_data[320],
                             in_data[205],
                             in_data[315]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [63:0] lut_273_table = 64'b0000000000000000111000001111000011110000111111001111010011111100;
    wire [5:0] lut_273_select = {
                             in_data[611],
                             in_data[257],
                             in_data[756],
                             in_data[187],
                             in_data[623],
                             in_data[284]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [63:0] lut_274_table = 64'b1111000011110000111101011111000000110000001100000011000000110000;
    wire [5:0] lut_274_select = {
                             in_data[329],
                             in_data[171],
                             in_data[64],
                             in_data[343],
                             in_data[130],
                             in_data[365]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [63:0] lut_275_table = 64'b0000001000001010001010101010101000000010001000100010101000101010;
    wire [5:0] lut_275_select = {
                             in_data[111],
                             in_data[713],
                             in_data[35],
                             in_data[631],
                             in_data[75],
                             in_data[154]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [63:0] lut_276_table = 64'b1010101110101111000010101010101010101011101011110000101010101010;
    wire [5:0] lut_276_select = {
                             in_data[224],
                             in_data[772],
                             in_data[78],
                             in_data[557],
                             in_data[751],
                             in_data[714]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [63:0] lut_277_table = 64'b0000000000000000000000000000000011001111110011111100110011001100;
    wire [5:0] lut_277_select = {
                             in_data[173],
                             in_data[292],
                             in_data[116],
                             in_data[501],
                             in_data[715],
                             in_data[31]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [63:0] lut_278_table = 64'b1111111100001010111111111010101011111111100010101111111110101010;
    wire [5:0] lut_278_select = {
                             in_data[310],
                             in_data[766],
                             in_data[102],
                             in_data[530],
                             in_data[534],
                             in_data[630]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [63:0] lut_279_table = 64'b1111110011111011110100001111100011111100111111111111100011111100;
    wire [5:0] lut_279_select = {
                             in_data[85],
                             in_data[709],
                             in_data[438],
                             in_data[434],
                             in_data[542],
                             in_data[95]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [63:0] lut_280_table = 64'b1111111111111111110101001101000011110001111100011111000101110001;
    wire [5:0] lut_280_select = {
                             in_data[182],
                             in_data[720],
                             in_data[90],
                             in_data[159],
                             in_data[323],
                             in_data[340]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [63:0] lut_281_table = 64'b0111001101110011001100100011001001110011011101110011000001110010;
    wire [5:0] lut_281_select = {
                             in_data[158],
                             in_data[215],
                             in_data[129],
                             in_data[276],
                             in_data[513],
                             in_data[314]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [63:0] lut_282_table = 64'b0000110000000000000000000000000011001100111111110000000000000000;
    wire [5:0] lut_282_select = {
                             in_data[305],
                             in_data[410],
                             in_data[127],
                             in_data[767],
                             in_data[551],
                             in_data[476]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [63:0] lut_283_table = 64'b1010101000001010111010100000000010101010000010001111101000000000;
    wire [5:0] lut_283_select = {
                             in_data[65],
                             in_data[321],
                             in_data[625],
                             in_data[175],
                             in_data[312],
                             in_data[570]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [63:0] lut_284_table = 64'b0001000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_284_select = {
                             in_data[356],
                             in_data[392],
                             in_data[658],
                             in_data[695],
                             in_data[169],
                             in_data[418]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [63:0] lut_285_table = 64'b1111111100110011111011100010001011111111001100111110111000110011;
    wire [5:0] lut_285_select = {
                             in_data[782],
                             in_data[443],
                             in_data[375],
                             in_data[477],
                             in_data[378],
                             in_data[298]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [63:0] lut_286_table = 64'b0000000000000000000011010000110100000000000001010000111100001111;
    wire [5:0] lut_286_select = {
                             in_data[219],
                             in_data[653],
                             in_data[81],
                             in_data[462],
                             in_data[497],
                             in_data[417]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [63:0] lut_287_table = 64'b0010000010110000101100001111000000000000000000000000000000110000;
    wire [5:0] lut_287_select = {
                             in_data[680],
                             in_data[638],
                             in_data[424],
                             in_data[377],
                             in_data[254],
                             in_data[708]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [63:0] lut_288_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_288_select = {
                             in_data[707],
                             in_data[283],
                             in_data[616],
                             in_data[579],
                             in_data[669],
                             in_data[316]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [63:0] lut_289_table = 64'b1111111101010101111111110000000011111111010101011111111100000000;
    wire [5:0] lut_289_select = {
                             in_data[190],
                             in_data[736],
                             in_data[133],
                             in_data[366],
                             in_data[391],
                             in_data[98]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [63:0] lut_290_table = 64'b1111111111101110111111111110111011111111111111111110111011101110;
    wire [5:0] lut_290_select = {
                             in_data[660],
                             in_data[155],
                             in_data[406],
                             in_data[3],
                             in_data[275],
                             in_data[201]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [63:0] lut_291_table = 64'b0000000000000000000000000000000000000000000000010000000000000011;
    wire [5:0] lut_291_select = {
                             in_data[577],
                             in_data[143],
                             in_data[496],
                             in_data[99],
                             in_data[231],
                             in_data[132]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [63:0] lut_292_table = 64'b0001000100000000000100000000000000010001000100010001000100010001;
    wire [5:0] lut_292_select = {
                             in_data[247],
                             in_data[337],
                             in_data[165],
                             in_data[141],
                             in_data[735],
                             in_data[711]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [63:0] lut_293_table = 64'b0000000000000000100000001000000011111111111111101111111111111111;
    wire [5:0] lut_293_select = {
                             in_data[516],
                             in_data[71],
                             in_data[53],
                             in_data[505],
                             in_data[307],
                             in_data[774]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [63:0] lut_294_table = 64'b0101010101010101010101010101010101010000010101010101000001010101;
    wire [5:0] lut_294_select = {
                             in_data[397],
                             in_data[543],
                             in_data[522],
                             in_data[635],
                             in_data[672],
                             in_data[273]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [63:0] lut_295_table = 64'b0000000011110000000000000000000011110000111111111111000011111111;
    wire [5:0] lut_295_select = {
                             in_data[467],
                             in_data[637],
                             in_data[608],
                             in_data[260],
                             in_data[194],
                             in_data[704]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [63:0] lut_296_table = 64'b0011001100110001011101110011001100110011000100010111011100110001;
    wire [5:0] lut_296_select = {
                             in_data[644],
                             in_data[341],
                             in_data[678],
                             in_data[289],
                             in_data[269],
                             in_data[429]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [63:0] lut_297_table = 64'b1101101100001011110111110000111111001011000010111101111100001111;
    wire [5:0] lut_297_select = {
                             in_data[309],
                             in_data[91],
                             in_data[367],
                             in_data[350],
                             in_data[547],
                             in_data[629]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [63:0] lut_298_table = 64'b1111111111111100111111111100110011111111111111001111111111001100;
    wire [5:0] lut_298_select = {
                             in_data[393],
                             in_data[56],
                             in_data[622],
                             in_data[436],
                             in_data[294],
                             in_data[639]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [63:0] lut_299_table = 64'b1110101011101010101010101010101011101110111010101010101010101010;
    wire [5:0] lut_299_select = {
                             in_data[673],
                             in_data[262],
                             in_data[728],
                             in_data[279],
                             in_data[521],
                             in_data[352]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [63:0] lut_300_table = 64'b0000000000000000000000000000000000110011000100110000001100000011;
    wire [5:0] lut_300_select = {
                             in_data[131],
                             in_data[399],
                             in_data[757],
                             in_data[665],
                             in_data[583],
                             in_data[750]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [63:0] lut_301_table = 64'b1111001111110011111100111111001111110011111100111111001111110011;
    wire [5:0] lut_301_select = {
                             in_data[390],
                             in_data[22],
                             in_data[243],
                             in_data[191],
                             in_data[490],
                             in_data[72]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [63:0] lut_302_table = 64'b1111111111111110111101110000000011111111011111111111111100000000;
    wire [5:0] lut_302_select = {
                             in_data[134],
                             in_data[396],
                             in_data[491],
                             in_data[318],
                             in_data[40],
                             in_data[363]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [63:0] lut_303_table = 64'b1110111111001111110011001100110011111111111011111100110011001100;
    wire [5:0] lut_303_select = {
                             in_data[761],
                             in_data[370],
                             in_data[688],
                             in_data[607],
                             in_data[234],
                             in_data[29]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [63:0] lut_304_table = 64'b1111001111110011001100110011001111100101110001010010001010100011;
    wire [5:0] lut_304_select = {
                             in_data[572],
                             in_data[302],
                             in_data[96],
                             in_data[416],
                             in_data[242],
                             in_data[357]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [63:0] lut_305_table = 64'b0000000000000000000000000000000000000000111111110000000001110101;
    wire [5:0] lut_305_select = {
                             in_data[682],
                             in_data[667],
                             in_data[189],
                             in_data[643],
                             in_data[666],
                             in_data[465]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [63:0] lut_306_table = 64'b0000000000000000001000000000000001010101010101010101010101010101;
    wire [5:0] lut_306_select = {
                             in_data[237],
                             in_data[89],
                             in_data[278],
                             in_data[506],
                             in_data[771],
                             in_data[209]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [63:0] lut_307_table = 64'b0000000000000000000000000101000000000000000000000000000001010000;
    wire [5:0] lut_307_select = {
                             in_data[452],
                             in_data[536],
                             in_data[676],
                             in_data[431],
                             in_data[777],
                             in_data[555]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [63:0] lut_308_table = 64'b1011001100110011001000100010001000111011001100110011001100110011;
    wire [5:0] lut_308_select = {
                             in_data[217],
                             in_data[358],
                             in_data[446],
                             in_data[562],
                             in_data[270],
                             in_data[123]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [63:0] lut_309_table = 64'b1010000011111010111110101111111100000000101000001010000010100000;
    wire [5:0] lut_309_select = {
                             in_data[409],
                             in_data[207],
                             in_data[287],
                             in_data[227],
                             in_data[114],
                             in_data[239]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [63:0] lut_310_table = 64'b1100111111111111110011001100110011111111111111111100110011001101;
    wire [5:0] lut_310_select = {
                             in_data[722],
                             in_data[193],
                             in_data[208],
                             in_data[42],
                             in_data[691],
                             in_data[422]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [63:0] lut_311_table = 64'b0011101111111111000100011101111110111111111011110000100011001100;
    wire [5:0] lut_311_select = {
                             in_data[651],
                             in_data[268],
                             in_data[685],
                             in_data[746],
                             in_data[566],
                             in_data[440]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [63:0] lut_312_table = 64'b0100000011110000010000001111000000000000010100000000000001010000;
    wire [5:0] lut_312_select = {
                             in_data[360],
                             in_data[336],
                             in_data[101],
                             in_data[656],
                             in_data[780],
                             in_data[94]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [63:0] lut_313_table = 64'b1111111111111111111111111111111110110010101100101111001011110010;
    wire [5:0] lut_313_select = {
                             in_data[453],
                             in_data[558],
                             in_data[252],
                             in_data[385],
                             in_data[546],
                             in_data[76]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [63:0] lut_314_table = 64'b1011101010111010111110111011101010111011101110111111101110111010;
    wire [5:0] lut_314_select = {
                             in_data[504],
                             in_data[726],
                             in_data[66],
                             in_data[172],
                             in_data[550],
                             in_data[510]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [63:0] lut_315_table = 64'b1111111111111101010101010101010111111111111111110101010101010101;
    wire [5:0] lut_315_select = {
                             in_data[773],
                             in_data[621],
                             in_data[586],
                             in_data[69],
                             in_data[282],
                             in_data[265]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [63:0] lut_316_table = 64'b1111010111110000111111101110101011110101111100001111000010101010;
    wire [5:0] lut_316_select = {
                             in_data[734],
                             in_data[156],
                             in_data[299],
                             in_data[486],
                             in_data[118],
                             in_data[326]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [63:0] lut_317_table = 64'b0000010100000101000001010000010100000101000001010000010100000101;
    wire [5:0] lut_317_select = {
                             in_data[142],
                             in_data[88],
                             in_data[383],
                             in_data[333],
                             in_data[748],
                             in_data[604]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [63:0] lut_318_table = 64'b1111111100000000111111110000000011111111111111111111111111111111;
    wire [5:0] lut_318_select = {
                             in_data[571],
                             in_data[744],
                             in_data[548],
                             in_data[697],
                             in_data[618],
                             in_data[703]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [63:0] lut_319_table = 64'b0000000000000000111110110000001100000000000000001111001100000000;
    wire [5:0] lut_319_select = {
                             in_data[12],
                             in_data[508],
                             in_data[574],
                             in_data[692],
                             in_data[747],
                             in_data[11]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [63:0] lut_320_table = 64'b1100110011001100000000000000000011001100110010001100110111011101;
    wire [5:0] lut_320_select = {
                             in_data[567],
                             in_data[553],
                             in_data[32],
                             in_data[110],
                             in_data[355],
                             in_data[166]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [63:0] lut_321_table = 64'b0000000000000000010001000000010000000000000000001100110111001101;
    wire [5:0] lut_321_select = {
                             in_data[176],
                             in_data[180],
                             in_data[528],
                             in_data[663],
                             in_data[624],
                             in_data[92]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [63:0] lut_322_table = 64'b1111111111111111111100001111000011111111111111111111111111111000;
    wire [5:0] lut_322_select = {
                             in_data[345],
                             in_data[414],
                             in_data[471],
                             in_data[151],
                             in_data[285],
                             in_data[25]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [63:0] lut_323_table = 64'b0000000011111011000000001111001100000000111100000000000011110000;
    wire [5:0] lut_323_select = {
                             in_data[466],
                             in_data[485],
                             in_data[342],
                             in_data[233],
                             in_data[334],
                             in_data[687]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [63:0] lut_324_table = 64'b1101111111001110111111111100111011011100111011101101110011111110;
    wire [5:0] lut_324_select = {
                             in_data[328],
                             in_data[413],
                             in_data[186],
                             in_data[210],
                             in_data[584],
                             in_data[293]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [63:0] lut_325_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_325_select = {
                             in_data[753],
                             in_data[313],
                             in_data[384],
                             in_data[645],
                             in_data[731],
                             in_data[614]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [63:0] lut_326_table = 64'b1111111011101110111111111110111011101110101010101110101010101010;
    wire [5:0] lut_326_select = {
                             in_data[769],
                             in_data[82],
                             in_data[41],
                             in_data[23],
                             in_data[218],
                             in_data[236]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [63:0] lut_327_table = 64'b0000000000000000000000000000000000000011000000110000001100000011;
    wire [5:0] lut_327_select = {
                             in_data[640],
                             in_data[14],
                             in_data[420],
                             in_data[192],
                             in_data[484],
                             in_data[9]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [63:0] lut_328_table = 64'b1111111110101010111111111010101011111111101010101111111110101010;
    wire [5:0] lut_328_select = {
                             in_data[526],
                             in_data[671],
                             in_data[124],
                             in_data[447],
                             in_data[759],
                             in_data[93]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [63:0] lut_329_table = 64'b1111010011100100111111111111111100000000000000000100010001000100;
    wire [5:0] lut_329_select = {
                             in_data[382],
                             in_data[261],
                             in_data[195],
                             in_data[13],
                             in_data[179],
                             in_data[712]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [63:0] lut_330_table = 64'b0000000001000101011100000111011100000000010101010111000001110111;
    wire [5:0] lut_330_select = {
                             in_data[106],
                             in_data[455],
                             in_data[601],
                             in_data[147],
                             in_data[509],
                             in_data[520]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [63:0] lut_331_table = 64'b1010001000000000111110111111000011111111110010001111111111111000;
    wire [5:0] lut_331_select = {
                             in_data[636],
                             in_data[605],
                             in_data[439],
                             in_data[444],
                             in_data[398],
                             in_data[525]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [63:0] lut_332_table = 64'b1111111111111100111111001100000011111111111111111111111111111100;
    wire [5:0] lut_332_select = {
                             in_data[719],
                             in_data[74],
                             in_data[73],
                             in_data[609],
                             in_data[595],
                             in_data[450]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [63:0] lut_333_table = 64'b0010000010100000101010101010101010100000101000001111101111111011;
    wire [5:0] lut_333_select = {
                             in_data[259],
                             in_data[122],
                             in_data[778],
                             in_data[369],
                             in_data[776],
                             in_data[146]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [63:0] lut_334_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_334_select = {
                             in_data[353],
                             in_data[34],
                             in_data[701],
                             in_data[113],
                             in_data[26],
                             in_data[538]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [63:0] lut_335_table = 64'b0000000000000000110011000000000011001100010000001100110011001100;
    wire [5:0] lut_335_select = {
                             in_data[655],
                             in_data[330],
                             in_data[620],
                             in_data[63],
                             in_data[544],
                             in_data[308]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [63:0] lut_336_table = 64'b1111011011111111111111111111111111111110111111101111111011111110;
    wire [5:0] lut_336_select = {
                             in_data[433],
                             in_data[763],
                             in_data[738],
                             in_data[304],
                             in_data[593],
                             in_data[153]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [63:0] lut_337_table = 64'b1110111111001111111111111111111110101010100011101010111010101110;
    wire [5:0] lut_337_select = {
                             in_data[626],
                             in_data[432],
                             in_data[17],
                             in_data[411],
                             in_data[44],
                             in_data[202]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [63:0] lut_338_table = 64'b1111111111111111101110011000100011111111110111011101110111011101;
    wire [5:0] lut_338_select = {
                             in_data[684],
                             in_data[181],
                             in_data[535],
                             in_data[38],
                             in_data[598],
                             in_data[325]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [63:0] lut_339_table = 64'b1010101000000000111111111010101010101010000000001111111110101010;
    wire [5:0] lut_339_select = {
                             in_data[137],
                             in_data[650],
                             in_data[599],
                             in_data[589],
                             in_data[770],
                             in_data[511]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [63:0] lut_340_table = 64'b1010101010101010111111111110111010101010000000000000000001010101;
    wire [5:0] lut_340_select = {
                             in_data[628],
                             in_data[649],
                             in_data[664],
                             in_data[752],
                             in_data[395],
                             in_data[633]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [63:0] lut_341_table = 64'b1000000010000000111001000000010010000100100001001110010010100101;
    wire [5:0] lut_341_select = {
                             in_data[250],
                             in_data[160],
                             in_data[472],
                             in_data[515],
                             in_data[573],
                             in_data[578]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [63:0] lut_342_table = 64'b0110011000100000001000100010000001110111011101110010001000100011;
    wire [5:0] lut_342_select = {
                             in_data[152],
                             in_data[373],
                             in_data[603],
                             in_data[721],
                             in_data[606],
                             in_data[463]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [63:0] lut_343_table = 64'b1111111111111111111111111111111100000000000000000101010101010100;
    wire [5:0] lut_343_select = {
                             in_data[499],
                             in_data[662],
                             in_data[754],
                             in_data[419],
                             in_data[500],
                             in_data[563]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [63:0] lut_344_table = 64'b1111110011111100110011001100110011111100111111001100110011001100;
    wire [5:0] lut_344_select = {
                             in_data[232],
                             in_data[575],
                             in_data[51],
                             in_data[407],
                             in_data[518],
                             in_data[762]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [63:0] lut_345_table = 64'b0011000100110001001100010011000100110001001100110011001100110011;
    wire [5:0] lut_345_select = {
                             in_data[613],
                             in_data[706],
                             in_data[112],
                             in_data[311],
                             in_data[430],
                             in_data[693]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [63:0] lut_346_table = 64'b0000000000000000000000000000000011110000111100001111110111111101;
    wire [5:0] lut_346_select = {
                             in_data[681],
                             in_data[482],
                             in_data[699],
                             in_data[495],
                             in_data[612],
                             in_data[581]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [63:0] lut_347_table = 64'b1010000010101010101100001111101000000000101010100000000011101110;
    wire [5:0] lut_347_select = {
                             in_data[381],
                             in_data[46],
                             in_data[322],
                             in_data[460],
                             in_data[729],
                             in_data[657]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [63:0] lut_348_table = 64'b0000000000000000001000000010001000000000000000000011001100110011;
    wire [5:0] lut_348_select = {
                             in_data[675],
                             in_data[203],
                             in_data[20],
                             in_data[62],
                             in_data[229],
                             in_data[674]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [63:0] lut_349_table = 64'b0011001100110011000000000000000011111111111111110010000010110011;
    wire [5:0] lut_349_select = {
                             in_data[677],
                             in_data[512],
                             in_data[324],
                             in_data[37],
                             in_data[412],
                             in_data[481]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [63:0] lut_350_table = 64'b0001000100000001000100010000000100010001000000010001000100000001;
    wire [5:0] lut_350_select = {
                             in_data[255],
                             in_data[61],
                             in_data[545],
                             in_data[461],
                             in_data[277],
                             in_data[221]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [63:0] lut_351_table = 64'b1111000011111010111100001111101011110000111110101111000011111010;
    wire [5:0] lut_351_select = {
                             in_data[591],
                             in_data[19],
                             in_data[387],
                             in_data[349],
                             in_data[1],
                             in_data[351]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [63:0] lut_352_table = 64'b1000000011110000000000001111000011110000111111011111000011111010;
    wire [5:0] lut_352_select = {
                             in_data[178],
                             in_data[28],
                             in_data[368],
                             in_data[300],
                             in_data[139],
                             in_data[80]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [63:0] lut_353_table = 64'b0101111101010111000101010000010101011111000001010001011100000101;
    wire [5:0] lut_353_select = {
                             in_data[272],
                             in_data[402],
                             in_data[710],
                             in_data[540],
                             in_data[128],
                             in_data[264]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [63:0] lut_354_table = 64'b0000111100001111100011111111111100001111000011110000111110001111;
    wire [5:0] lut_354_select = {
                             in_data[281],
                             in_data[241],
                             in_data[258],
                             in_data[266],
                             in_data[196],
                             in_data[52]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [63:0] lut_355_table = 64'b0111000001110000000000000000000011110011111100110000000000000000;
    wire [5:0] lut_355_select = {
                             in_data[145],
                             in_data[290],
                             in_data[5],
                             in_data[428],
                             in_data[537],
                             in_data[492]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [63:0] lut_356_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_356_select = {
                             in_data[119],
                             in_data[404],
                             in_data[223],
                             in_data[27],
                             in_data[6],
                             in_data[117]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [63:0] lut_357_table = 64'b1111111111001101111111111100110001000000110011000000000011001100;
    wire [5:0] lut_357_select = {
                             in_data[523],
                             in_data[83],
                             in_data[457],
                             in_data[58],
                             in_data[376],
                             in_data[253]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [63:0] lut_358_table = 64'b1111111111111111111111111111111111111111111111111110111100000000;
    wire [5:0] lut_358_select = {
                             in_data[163],
                             in_data[554],
                             in_data[109],
                             in_data[7],
                             in_data[531],
                             in_data[449]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [63:0] lut_359_table = 64'b0101110101000100000000000000000011111111111111111101110001000101;
    wire [5:0] lut_359_select = {
                             in_data[339],
                             in_data[48],
                             in_data[54],
                             in_data[617],
                             in_data[646],
                             in_data[86]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [63:0] lut_360_table = 64'b1111111111111111000001000000000011111111111111111111111011111111;
    wire [5:0] lut_360_select = {
                             in_data[517],
                             in_data[425],
                             in_data[458],
                             in_data[36],
                             in_data[775],
                             in_data[696]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [63:0] lut_361_table = 64'b0101010101010101000000000000000001010101010101010101010101010101;
    wire [5:0] lut_361_select = {
                             in_data[427],
                             in_data[585],
                             in_data[50],
                             in_data[779],
                             in_data[724],
                             in_data[582]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [63:0] lut_362_table = 64'b0001000100010001000000000000000001010111010101110000000000000000;
    wire [5:0] lut_362_select = {
                             in_data[451],
                             in_data[317],
                             in_data[228],
                             in_data[435],
                             in_data[718],
                             in_data[256]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [63:0] lut_363_table = 64'b1111111111111111111111111111111110101111001011001010111100101100;
    wire [5:0] lut_363_select = {
                             in_data[442],
                             in_data[115],
                             in_data[415],
                             in_data[214],
                             in_data[246],
                             in_data[204]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [63:0] lut_364_table = 64'b1010101110101011101010101010101100001010000010100000101000001010;
    wire [5:0] lut_364_select = {
                             in_data[488],
                             in_data[619],
                             in_data[338],
                             in_data[332],
                             in_data[388],
                             in_data[379]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [63:0] lut_365_table = 64'b1010111110101111101011111010111100001111000011110000111100001111;
    wire [5:0] lut_365_select = {
                             in_data[743],
                             in_data[104],
                             in_data[138],
                             in_data[372],
                             in_data[170],
                             in_data[354]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [63:0] lut_366_table = 64'b1111111111111111111101111111000111111111111101011111010101110000;
    wire [5:0] lut_366_select = {
                             in_data[77],
                             in_data[105],
                             in_data[198],
                             in_data[67],
                             in_data[723],
                             in_data[647]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [63:0] lut_367_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_367_select = {
                             in_data[288],
                             in_data[21],
                             in_data[527],
                             in_data[760],
                             in_data[594],
                             in_data[197]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [63:0] lut_368_table = 64'b0101010101010101010101010101111101000100010101010101010101010101;
    wire [5:0] lut_368_select = {
                             in_data[100],
                             in_data[749],
                             in_data[319],
                             in_data[49],
                             in_data[725],
                             in_data[296]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [63:0] lut_369_table = 64'b1111111111111111111111111111111111111111010101011111111100000000;
    wire [5:0] lut_369_select = {
                             in_data[426],
                             in_data[251],
                             in_data[745],
                             in_data[700],
                             in_data[758],
                             in_data[167]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [63:0] lut_370_table = 64'b1111011111110000000000000011000011110111111100000010000000100000;
    wire [5:0] lut_370_select = {
                             in_data[560],
                             in_data[271],
                             in_data[654],
                             in_data[549],
                             in_data[741],
                             in_data[519]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [63:0] lut_371_table = 64'b1101010111011101010101011101010111011101110111011101110111011101;
    wire [5:0] lut_371_select = {
                             in_data[740],
                             in_data[68],
                             in_data[361],
                             in_data[199],
                             in_data[580],
                             in_data[213]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [63:0] lut_372_table = 64'b1110111010001110111111111111111111001110100011101110111011101111;
    wire [5:0] lut_372_select = {
                             in_data[474],
                             in_data[183],
                             in_data[648],
                             in_data[344],
                             in_data[157],
                             in_data[177]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [63:0] lut_373_table = 64'b1111111111111111111111111111111111000000111100001111000011110000;
    wire [5:0] lut_373_select = {
                             in_data[689],
                             in_data[507],
                             in_data[742],
                             in_data[539],
                             in_data[10],
                             in_data[374]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [63:0] lut_374_table = 64'b0111001100000000111100111111000101000000111100001111000011110000;
    wire [5:0] lut_374_select = {
                             in_data[524],
                             in_data[362],
                             in_data[454],
                             in_data[348],
                             in_data[576],
                             in_data[18]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [63:0] lut_375_table = 64'b0001000000010000001100010111000111111011111100110011001100110011;
    wire [5:0] lut_375_select = {
                             in_data[371],
                             in_data[263],
                             in_data[136],
                             in_data[274],
                             in_data[347],
                             in_data[470]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [63:0] lut_376_table = 64'b1111111111110011111111111111001111111111111100111111111111110011;
    wire [5:0] lut_376_select = {
                             in_data[249],
                             in_data[561],
                             in_data[248],
                             in_data[456],
                             in_data[627],
                             in_data[225]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [63:0] lut_377_table = 64'b1111101011111111101010101111111111111010111111111010101011111111;
    wire [5:0] lut_377_select = {
                             in_data[15],
                             in_data[364],
                             in_data[212],
                             in_data[331],
                             in_data[55],
                             in_data[135]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [63:0] lut_378_table = 64'b1111111111111111000011111010111111111111111111110000101010001111;
    wire [5:0] lut_378_select = {
                             in_data[502],
                             in_data[565],
                             in_data[401],
                             in_data[188],
                             in_data[335],
                             in_data[498]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [63:0] lut_379_table = 64'b1111111111111111111111111100110011001111110011101100110011001100;
    wire [5:0] lut_379_select = {
                             in_data[514],
                             in_data[634],
                             in_data[683],
                             in_data[162],
                             in_data[405],
                             in_data[559]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [63:0] lut_380_table = 64'b1111111111111111111111111111111111111111111111111111100011111000;
    wire [5:0] lut_380_select = {
                             in_data[120],
                             in_data[610],
                             in_data[478],
                             in_data[97],
                             in_data[185],
                             in_data[327]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [63:0] lut_381_table = 64'b0000000000000000000000001100110011001100111111111100110011111111;
    wire [5:0] lut_381_select = {
                             in_data[400],
                             in_data[24],
                             in_data[483],
                             in_data[33],
                             in_data[489],
                             in_data[702]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [63:0] lut_382_table = 64'b0101010101010101010101011101110100000000000000000000000000000000;
    wire [5:0] lut_382_select = {
                             in_data[238],
                             in_data[533],
                             in_data[698],
                             in_data[493],
                             in_data[4],
                             in_data[216]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [63:0] lut_383_table = 64'b1111111111111101110000000000000011111111111111111010100010000000;
    wire [5:0] lut_383_select = {
                             in_data[568],
                             in_data[494],
                             in_data[448],
                             in_data[389],
                             in_data[39],
                             in_data[244]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [63:0] lut_384_table = 64'b1111111111110001111111110111000111111111111100001111111101110010;
    wire [5:0] lut_384_select = {
                             in_data[730],
                             in_data[30],
                             in_data[564],
                             in_data[148],
                             in_data[301],
                             in_data[0]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [63:0] lut_385_table = 64'b0000000000000000000000000000000011111111111111111111111100000000;
    wire [5:0] lut_385_select = {
                             in_data[226],
                             in_data[764],
                             in_data[149],
                             in_data[783],
                             in_data[781],
                             in_data[140]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [63:0] lut_386_table = 64'b1111111100110011111111110011001111111111001100111111111100110011;
    wire [5:0] lut_386_select = {
                             in_data[670],
                             in_data[359],
                             in_data[480],
                             in_data[280],
                             in_data[403],
                             in_data[768]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [63:0] lut_387_table = 64'b1100000011000000000000000000000011111101111111110100110101001101;
    wire [5:0] lut_387_select = {
                             in_data[386],
                             in_data[184],
                             in_data[84],
                             in_data[245],
                             in_data[200],
                             in_data[739]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [63:0] lut_388_table = 64'b1111111111111110111111111111111111111111000000001111111100000000;
    wire [5:0] lut_388_select = {
                             in_data[468],
                             in_data[2],
                             in_data[211],
                             in_data[755],
                             in_data[732],
                             in_data[108]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [63:0] lut_389_table = 64'b0000000000010001000000000001000100000000000100010000000000010001;
    wire [5:0] lut_389_select = {
                             in_data[716],
                             in_data[590],
                             in_data[592],
                             in_data[394],
                             in_data[206],
                             in_data[174]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [63:0] lut_390_table = 64'b1111111111111111111111111111111100000000000101010000000000010000;
    wire [5:0] lut_390_select = {
                             in_data[634],
                             in_data[781],
                             in_data[437],
                             in_data[60],
                             in_data[475],
                             in_data[445]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [63:0] lut_391_table = 64'b1010111110101111101011111010111111111111111011111010111110101111;
    wire [5:0] lut_391_select = {
                             in_data[518],
                             in_data[356],
                             in_data[0],
                             in_data[316],
                             in_data[21],
                             in_data[284]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [63:0] lut_392_table = 64'b1111000011110000111100001111000011110000111100011111000011110000;
    wire [5:0] lut_392_select = {
                             in_data[278],
                             in_data[45],
                             in_data[33],
                             in_data[595],
                             in_data[366],
                             in_data[552]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [63:0] lut_393_table = 64'b0000111110001111100011111000111100001111000011110000111100001111;
    wire [5:0] lut_393_select = {
                             in_data[590],
                             in_data[701],
                             in_data[5],
                             in_data[180],
                             in_data[714],
                             in_data[560]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [63:0] lut_394_table = 64'b1000111110101111101011111010111111110000111110101111101011111010;
    wire [5:0] lut_394_select = {
                             in_data[288],
                             in_data[503],
                             in_data[530],
                             in_data[359],
                             in_data[112],
                             in_data[734]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [63:0] lut_395_table = 64'b1111111100110011111111110011001111111111001100111111111100110011;
    wire [5:0] lut_395_select = {
                             in_data[721],
                             in_data[227],
                             in_data[512],
                             in_data[588],
                             in_data[543],
                             in_data[674]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [63:0] lut_396_table = 64'b1111111100001111111111110000000111111111000011111111111100000101;
    wire [5:0] lut_396_select = {
                             in_data[140],
                             in_data[103],
                             in_data[155],
                             in_data[237],
                             in_data[171],
                             in_data[174]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [63:0] lut_397_table = 64'b1111111111111111111111111111111101010000010100000000000000001000;
    wire [5:0] lut_397_select = {
                             in_data[344],
                             in_data[347],
                             in_data[447],
                             in_data[461],
                             in_data[28],
                             in_data[91]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [63:0] lut_398_table = 64'b1111111111110101111111110101010011111111111101111111111111110111;
    wire [5:0] lut_398_select = {
                             in_data[492],
                             in_data[746],
                             in_data[651],
                             in_data[220],
                             in_data[282],
                             in_data[352]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [63:0] lut_399_table = 64'b1111111111111111111111001111111001011111111111111110111011111110;
    wire [5:0] lut_399_select = {
                             in_data[520],
                             in_data[272],
                             in_data[259],
                             in_data[686],
                             in_data[738],
                             in_data[273]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [63:0] lut_400_table = 64'b0000111100001111000011110000111111111111000011111111111100001111;
    wire [5:0] lut_400_select = {
                             in_data[717],
                             in_data[42],
                             in_data[453],
                             in_data[185],
                             in_data[10],
                             in_data[110]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [63:0] lut_401_table = 64'b0000000000000000000000000111011100000000000000000000000000010001;
    wire [5:0] lut_401_select = {
                             in_data[154],
                             in_data[657],
                             in_data[631],
                             in_data[113],
                             in_data[331],
                             in_data[228]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [63:0] lut_402_table = 64'b1010101111111111000000000000000011111111111111110000010101010111;
    wire [5:0] lut_402_select = {
                             in_data[574],
                             in_data[609],
                             in_data[187],
                             in_data[770],
                             in_data[51],
                             in_data[204]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [63:0] lut_403_table = 64'b0000000011110000000000001100000011110000111111111111000011111111;
    wire [5:0] lut_403_select = {
                             in_data[209],
                             in_data[41],
                             in_data[747],
                             in_data[441],
                             in_data[765],
                             in_data[478]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [63:0] lut_404_table = 64'b1011101100000000101110110000000011111111111111111111111111111111;
    wire [5:0] lut_404_select = {
                             in_data[371],
                             in_data[16],
                             in_data[567],
                             in_data[731],
                             in_data[539],
                             in_data[100]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [63:0] lut_405_table = 64'b0000111100001111000011110000111100001111000011110000111100001111;
    wire [5:0] lut_405_select = {
                             in_data[732],
                             in_data[604],
                             in_data[446],
                             in_data[568],
                             in_data[368],
                             in_data[696]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [63:0] lut_406_table = 64'b1010101010101010101010101010101011101010101010101010101010101010;
    wire [5:0] lut_406_select = {
                             in_data[58],
                             in_data[689],
                             in_data[725],
                             in_data[691],
                             in_data[349],
                             in_data[654]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [63:0] lut_407_table = 64'b1111111111111111110011001100110011111111111111111110110011001100;
    wire [5:0] lut_407_select = {
                             in_data[418],
                             in_data[666],
                             in_data[728],
                             in_data[15],
                             in_data[358],
                             in_data[53]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [63:0] lut_408_table = 64'b0000000000000000111100001111000000000000000000001100000011100000;
    wire [5:0] lut_408_select = {
                             in_data[381],
                             in_data[501],
                             in_data[306],
                             in_data[429],
                             in_data[274],
                             in_data[671]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [63:0] lut_409_table = 64'b0101000000000000111101010000000001010000101011011101010111111111;
    wire [5:0] lut_409_select = {
                             in_data[542],
                             in_data[678],
                             in_data[493],
                             in_data[267],
                             in_data[223],
                             in_data[462]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [63:0] lut_410_table = 64'b0000000000000000101010100000000011111111111111111011111110101010;
    wire [5:0] lut_410_select = {
                             in_data[291],
                             in_data[287],
                             in_data[385],
                             in_data[771],
                             in_data[777],
                             in_data[383]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [63:0] lut_411_table = 64'b0000000000000000111100001111111100000000000000001111000011110000;
    wire [5:0] lut_411_select = {
                             in_data[338],
                             in_data[162],
                             in_data[555],
                             in_data[242],
                             in_data[225],
                             in_data[29]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [63:0] lut_412_table = 64'b0000000000000000000000000001000000010000001100000011000001110001;
    wire [5:0] lut_412_select = {
                             in_data[334],
                             in_data[415],
                             in_data[136],
                             in_data[144],
                             in_data[135],
                             in_data[69]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [63:0] lut_413_table = 64'b1010101010101010111010101010101011101110111011101111111111101111;
    wire [5:0] lut_413_select = {
                             in_data[217],
                             in_data[733],
                             in_data[7],
                             in_data[336],
                             in_data[40],
                             in_data[362]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [63:0] lut_414_table = 64'b1100110001001100111111111101111101001100000000001111111111001100;
    wire [5:0] lut_414_select = {
                             in_data[584],
                             in_data[427],
                             in_data[193],
                             in_data[759],
                             in_data[212],
                             in_data[663]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [63:0] lut_415_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_415_select = {
                             in_data[55],
                             in_data[684],
                             in_data[495],
                             in_data[54],
                             in_data[6],
                             in_data[249]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [63:0] lut_416_table = 64'b1111001111110011111100111111001100110011111100000011001011110000;
    wire [5:0] lut_416_select = {
                             in_data[471],
                             in_data[64],
                             in_data[467],
                             in_data[457],
                             in_data[326],
                             in_data[36]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [63:0] lut_417_table = 64'b1111111110101011111111111010111111111111101011111011111100001111;
    wire [5:0] lut_417_select = {
                             in_data[121],
                             in_data[353],
                             in_data[425],
                             in_data[350],
                             in_data[750],
                             in_data[544]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [63:0] lut_418_table = 64'b0000101000001000000011110000101000001111000011110000111100001111;
    wire [5:0] lut_418_select = {
                             in_data[409],
                             in_data[585],
                             in_data[66],
                             in_data[498],
                             in_data[22],
                             in_data[693]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [63:0] lut_419_table = 64'b0111011101110111011101110101010111110101011101010111010101010101;
    wire [5:0] lut_419_select = {
                             in_data[569],
                             in_data[563],
                             in_data[258],
                             in_data[201],
                             in_data[687],
                             in_data[215]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [63:0] lut_420_table = 64'b0000001100100000000000110010000010101111101100111010111110110011;
    wire [5:0] lut_420_select = {
                             in_data[536],
                             in_data[198],
                             in_data[188],
                             in_data[608],
                             in_data[514],
                             in_data[147]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [63:0] lut_421_table = 64'b1100110000000000110011000000000011001100000000001101110101000101;
    wire [5:0] lut_421_select = {
                             in_data[145],
                             in_data[489],
                             in_data[294],
                             in_data[422],
                             in_data[321],
                             in_data[148]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [63:0] lut_422_table = 64'b1111111100010001111111110000000011111111000100011111111100000000;
    wire [5:0] lut_422_select = {
                             in_data[76],
                             in_data[405],
                             in_data[434],
                             in_data[618],
                             in_data[165],
                             in_data[395]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [63:0] lut_423_table = 64'b1111000111110111011100010000000111110001111101110111000100000001;
    wire [5:0] lut_423_select = {
                             in_data[531],
                             in_data[472],
                             in_data[301],
                             in_data[458],
                             in_data[256],
                             in_data[176]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [63:0] lut_424_table = 64'b0000000000000000000000000000000011011101110011000101010101000101;
    wire [5:0] lut_424_select = {
                             in_data[276],
                             in_data[236],
                             in_data[311],
                             in_data[77],
                             in_data[428],
                             in_data[160]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [63:0] lut_425_table = 64'b0000000000001000100010001110111000000000110011001100110011111111;
    wire [5:0] lut_425_select = {
                             in_data[516],
                             in_data[407],
                             in_data[715],
                             in_data[255],
                             in_data[443],
                             in_data[414]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [63:0] lut_426_table = 64'b1111111111110101011100010000000011111101110101010001000100000000;
    wire [5:0] lut_426_select = {
                             in_data[75],
                             in_data[372],
                             in_data[402],
                             in_data[742],
                             in_data[424],
                             in_data[124]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [63:0] lut_427_table = 64'b0000000000000000000100000001000000000000000000000101000001010000;
    wire [5:0] lut_427_select = {
                             in_data[80],
                             in_data[554],
                             in_data[111],
                             in_data[599],
                             in_data[707],
                             in_data[122]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [63:0] lut_428_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_428_select = {
                             in_data[169],
                             in_data[736],
                             in_data[292],
                             in_data[632],
                             in_data[783],
                             in_data[626]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [63:0] lut_429_table = 64'b1000000001110001000000000111000100000000010101010000000001010101;
    wire [5:0] lut_429_select = {
                             in_data[213],
                             in_data[35],
                             in_data[440],
                             in_data[581],
                             in_data[384],
                             in_data[150]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [63:0] lut_430_table = 64'b0010000000100000101110111011001100100010101000101111101111111111;
    wire [5:0] lut_430_select = {
                             in_data[720],
                             in_data[466],
                             in_data[751],
                             in_data[444],
                             in_data[183],
                             in_data[95]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [63:0] lut_431_table = 64'b0000110100001111000001000000111100001101000011110000010000001101;
    wire [5:0] lut_431_select = {
                             in_data[98],
                             in_data[591],
                             in_data[374],
                             in_data[191],
                             in_data[723],
                             in_data[309]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [63:0] lut_432_table = 64'b0000101000001010000010100000101010101111000011110000111100001111;
    wire [5:0] lut_432_select = {
                             in_data[342],
                             in_data[729],
                             in_data[647],
                             in_data[605],
                             in_data[59],
                             in_data[547]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [63:0] lut_433_table = 64'b0000000000000101000000000010111100000000000000000000111100001111;
    wire [5:0] lut_433_select = {
                             in_data[318],
                             in_data[580],
                             in_data[433],
                             in_data[635],
                             in_data[119],
                             in_data[583]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [63:0] lut_434_table = 64'b0000000011000100010001001100110000000000110011001100110011001100;
    wire [5:0] lut_434_select = {
                             in_data[206],
                             in_data[189],
                             in_data[650],
                             in_data[137],
                             in_data[577],
                             in_data[345]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [63:0] lut_435_table = 64'b0000000000000000111111001110100011101000101010001111111111111110;
    wire [5:0] lut_435_select = {
                             in_data[613],
                             in_data[640],
                             in_data[365],
                             in_data[172],
                             in_data[92],
                             in_data[194]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [63:0] lut_436_table = 64'b1111111111111111111111111111111111111010111110101111101011111010;
    wire [5:0] lut_436_select = {
                             in_data[315],
                             in_data[570],
                             in_data[252],
                             in_data[247],
                             in_data[11],
                             in_data[339]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [63:0] lut_437_table = 64'b1010111011111111000011100111111100000111000011110000000001001111;
    wire [5:0] lut_437_select = {
                             in_data[178],
                             in_data[628],
                             in_data[602],
                             in_data[411],
                             in_data[302],
                             in_data[578]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [63:0] lut_438_table = 64'b0101010001010100010000000100000011111111111111110000000000010000;
    wire [5:0] lut_438_select = {
                             in_data[261],
                             in_data[603],
                             in_data[62],
                             in_data[184],
                             in_data[233],
                             in_data[744]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [63:0] lut_439_table = 64'b1010000010100000101000001010000010100000101000001010000010100000;
    wire [5:0] lut_439_select = {
                             in_data[1],
                             in_data[50],
                             in_data[639],
                             in_data[438],
                             in_data[768],
                             in_data[576]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [63:0] lut_440_table = 64'b1111101100110000111111111111000000000000000000001111111111001100;
    wire [5:0] lut_440_select = {
                             in_data[549],
                             in_data[297],
                             in_data[523],
                             in_data[575],
                             in_data[661],
                             in_data[17]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [63:0] lut_441_table = 64'b1111111111111111110011001111111111101110111011101100010011101110;
    wire [5:0] lut_441_select = {
                             in_data[99],
                             in_data[665],
                             in_data[521],
                             in_data[699],
                             in_data[592],
                             in_data[323]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [63:0] lut_442_table = 64'b1010101011111111101010101010101010101010101011111010101010101010;
    wire [5:0] lut_442_select = {
                             in_data[329],
                             in_data[659],
                             in_data[545],
                             in_data[586],
                             in_data[34],
                             in_data[293]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [63:0] lut_443_table = 64'b0100010001000100010101010101010101000100010001000101010001000100;
    wire [5:0] lut_443_select = {
                             in_data[120],
                             in_data[151],
                             in_data[67],
                             in_data[44],
                             in_data[214],
                             in_data[566]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [63:0] lut_444_table = 64'b0000111100001100000011110000110100001111000011011000111100001111;
    wire [5:0] lut_444_select = {
                             in_data[504],
                             in_data[668],
                             in_data[515],
                             in_data[295],
                             in_data[27],
                             in_data[56]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [63:0] lut_445_table = 64'b0000000000000000000000001111111100000000111111110000000011111111;
    wire [5:0] lut_445_select = {
                             in_data[465],
                             in_data[662],
                             in_data[317],
                             in_data[506],
                             in_data[14],
                             in_data[389]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [63:0] lut_446_table = 64'b1111111111111111010100000101000011111111111111110101010101010101;
    wire [5:0] lut_446_select = {
                             in_data[403],
                             in_data[623],
                             in_data[745],
                             in_data[752],
                             in_data[420],
                             in_data[398]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [63:0] lut_447_table = 64'b1111111111111111111110101010000011111111111111111111111111111010;
    wire [5:0] lut_447_select = {
                             in_data[199],
                             in_data[128],
                             in_data[638],
                             in_data[219],
                             in_data[508],
                             in_data[431]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [63:0] lut_448_table = 64'b0000000000001100111011111100111100000000000000000000110011001101;
    wire [5:0] lut_448_select = {
                             in_data[529],
                             in_data[248],
                             in_data[179],
                             in_data[679],
                             in_data[129],
                             in_data[81]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [63:0] lut_449_table = 64'b0001110000000000000010000000110011110000111111111111000011111111;
    wire [5:0] lut_449_select = {
                             in_data[455],
                             in_data[63],
                             in_data[488],
                             in_data[540],
                             in_data[413],
                             in_data[669]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [63:0] lut_450_table = 64'b1111111100000000111111111011001011111111000000001111111100000000;
    wire [5:0] lut_450_select = {
                             in_data[268],
                             in_data[304],
                             in_data[97],
                             in_data[26],
                             in_data[724],
                             in_data[43]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [63:0] lut_451_table = 64'b0101000011011111010100001111111101010000110111110101000011011111;
    wire [5:0] lut_451_select = {
                             in_data[764],
                             in_data[727],
                             in_data[210],
                             in_data[386],
                             in_data[587],
                             in_data[460]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [63:0] lut_452_table = 64'b1111101011101010111111101110100010100000111110100100000011111110;
    wire [5:0] lut_452_select = {
                             in_data[468],
                             in_data[341],
                             in_data[553],
                             in_data[133],
                             in_data[325],
                             in_data[207]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [63:0] lut_453_table = 64'b1110111111101110111011111110111011101111111011101110111111101110;
    wire [5:0] lut_453_select = {
                             in_data[82],
                             in_data[704],
                             in_data[68],
                             in_data[483],
                             in_data[627],
                             in_data[528]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [63:0] lut_454_table = 64'b1100110011001100000011110000111111111100111111000010111100001111;
    wire [5:0] lut_454_select = {
                             in_data[675],
                             in_data[216],
                             in_data[226],
                             in_data[401],
                             in_data[633],
                             in_data[335]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [63:0] lut_455_table = 64'b0101010101011111000000000000010101010101010101010000000000000000;
    wire [5:0] lut_455_select = {
                             in_data[522],
                             in_data[509],
                             in_data[312],
                             in_data[367],
                             in_data[308],
                             in_data[396]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [63:0] lut_456_table = 64'b1111110011110000111111111111111111101100111000001111111111111111;
    wire [5:0] lut_456_select = {
                             in_data[83],
                             in_data[410],
                             in_data[619],
                             in_data[181],
                             in_data[582],
                             in_data[281]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [63:0] lut_457_table = 64'b0101010101010101010101011111111100000000000000000000000000010001;
    wire [5:0] lut_457_select = {
                             in_data[322],
                             in_data[454],
                             in_data[426],
                             in_data[23],
                             in_data[221],
                             in_data[146]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [63:0] lut_458_table = 64'b0000000000000000000000000000000000001100110011110000110011001111;
    wire [5:0] lut_458_select = {
                             in_data[388],
                             in_data[57],
                             in_data[125],
                             in_data[534],
                             in_data[749],
                             in_data[2]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [63:0] lut_459_table = 64'b0011001110111011001100111011001100110011101110110011001110110011;
    wire [5:0] lut_459_select = {
                             in_data[391],
                             in_data[104],
                             in_data[269],
                             in_data[557],
                             in_data[205],
                             in_data[361]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [63:0] lut_460_table = 64'b0000000001110000000000000000000011110000111111110101000011110000;
    wire [5:0] lut_460_select = {
                             in_data[442],
                             in_data[157],
                             in_data[369],
                             in_data[156],
                             in_data[8],
                             in_data[392]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [63:0] lut_461_table = 64'b1110110011111111111010001111111111101100111111111100100011101111;
    wire [5:0] lut_461_select = {
                             in_data[25],
                             in_data[115],
                             in_data[118],
                             in_data[589],
                             in_data[13],
                             in_data[562]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [63:0] lut_462_table = 64'b1111111111111111110011010100110011111111111111111100110101001100;
    wire [5:0] lut_462_select = {
                             in_data[307],
                             in_data[624],
                             in_data[319],
                             in_data[406],
                             in_data[480],
                             in_data[170]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [63:0] lut_463_table = 64'b0000000000110011000000000000000000110011001100110010000011111111;
    wire [5:0] lut_463_select = {
                             in_data[527],
                             in_data[132],
                             in_data[285],
                             in_data[251],
                             in_data[271],
                             in_data[450]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [63:0] lut_464_table = 64'b1111111111111111111111111111111111111111110011001111111111001100;
    wire [5:0] lut_464_select = {
                             in_data[629],
                             in_data[476],
                             in_data[298],
                             in_data[756],
                             in_data[594],
                             in_data[449]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [63:0] lut_465_table = 64'b0000111100001110000011110000111110101111000011111111111100001111;
    wire [5:0] lut_465_select = {
                             in_data[743],
                             in_data[253],
                             in_data[676],
                             in_data[484],
                             in_data[673],
                             in_data[46]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [63:0] lut_466_table = 64'b1111111110101010111111111010101011111111101110111111111110101011;
    wire [5:0] lut_466_select = {
                             in_data[463],
                             in_data[564],
                             in_data[257],
                             in_data[558],
                             in_data[517],
                             in_data[72]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [63:0] lut_467_table = 64'b1000111100001111000011110000110000001111000011110000111100001100;
    wire [5:0] lut_467_select = {
                             in_data[645],
                             in_data[737],
                             in_data[494],
                             in_data[93],
                             in_data[716],
                             in_data[741]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [63:0] lut_468_table = 64'b1111111101110111001100110011001111111111001100110011001100110011;
    wire [5:0] lut_468_select = {
                             in_data[740],
                             in_data[464],
                             in_data[203],
                             in_data[532],
                             in_data[290],
                             in_data[606]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [63:0] lut_469_table = 64'b0000000000001111000000000000000000000011001111110000001100000010;
    wire [5:0] lut_469_select = {
                             in_data[333],
                             in_data[435],
                             in_data[546],
                             in_data[652],
                             in_data[231],
                             in_data[755]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [63:0] lut_470_table = 64'b0000110000000000000011000000100011001111110011111100111111001111;
    wire [5:0] lut_470_select = {
                             in_data[234],
                             in_data[419],
                             in_data[763],
                             in_data[175],
                             in_data[131],
                             in_data[561]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [63:0] lut_471_table = 64'b0000000000000000000000001111111100000000000000000000000011111111;
    wire [5:0] lut_471_select = {
                             in_data[758],
                             in_data[351],
                             in_data[712],
                             in_data[706],
                             in_data[757],
                             in_data[238]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [63:0] lut_472_table = 64'b0000000000000000000011110000111100000000000000000000111100001111;
    wire [5:0] lut_472_select = {
                             in_data[642],
                             in_data[486],
                             in_data[102],
                             in_data[126],
                             in_data[664],
                             in_data[138]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [63:0] lut_473_table = 64'b1111111111111111010001000100010011111111111111111110110011001110;
    wire [5:0] lut_473_select = {
                             in_data[208],
                             in_data[596],
                             in_data[616],
                             in_data[116],
                             in_data[511],
                             in_data[346]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [63:0] lut_474_table = 64'b0000000000000000000000000000000000001111000011010000111100001111;
    wire [5:0] lut_474_select = {
                             in_data[481],
                             in_data[614],
                             in_data[718],
                             in_data[622],
                             in_data[767],
                             in_data[86]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [63:0] lut_475_table = 64'b0101010101010101110111010101010101010101010101010101010101010101;
    wire [5:0] lut_475_select = {
                             in_data[314],
                             in_data[108],
                             in_data[280],
                             in_data[142],
                             in_data[593],
                             in_data[513]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [63:0] lut_476_table = 64'b1111001100110001111100110011001101110011001100110011001100110011;
    wire [5:0] lut_476_select = {
                             in_data[762],
                             in_data[615],
                             in_data[601],
                             in_data[692],
                             in_data[377],
                             in_data[761]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [63:0] lut_477_table = 64'b0000000000000000000001010000010100000000000000000000110100000101;
    wire [5:0] lut_477_select = {
                             in_data[730],
                             in_data[130],
                             in_data[173],
                             in_data[360],
                             in_data[690],
                             in_data[357]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [63:0] lut_478_table = 64'b1111111111111111111111111111111111111111111111110000000011001110;
    wire [5:0] lut_478_select = {
                             in_data[680],
                             in_data[695],
                             in_data[697],
                             in_data[12],
                             in_data[65],
                             in_data[196]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [63:0] lut_479_table = 64'b1111111010111011111111110011001011111110111100111111111100100010;
    wire [5:0] lut_479_select = {
                             in_data[393],
                             in_data[327],
                             in_data[330],
                             in_data[773],
                             in_data[134],
                             in_data[775]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [63:0] lut_480_table = 64'b0000000000000000000000000000000000000000000000001111111111111111;
    wire [5:0] lut_480_select = {
                             in_data[182],
                             in_data[222],
                             in_data[143],
                             in_data[753],
                             in_data[19],
                             in_data[477]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [63:0] lut_481_table = 64'b0011001100110011001100110011001100010000001100110011001000110011;
    wire [5:0] lut_481_select = {
                             in_data[343],
                             in_data[735],
                             in_data[766],
                             in_data[32],
                             in_data[470],
                             in_data[778]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [63:0] lut_482_table = 64'b1111111111111111111110001111111011111110111111111110100011111000;
    wire [5:0] lut_482_select = {
                             in_data[535],
                             in_data[262],
                             in_data[340],
                             in_data[439],
                             in_data[620],
                             in_data[682]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [63:0] lut_483_table = 64'b1111011100110001111111110011000100010101000100010001010100010001;
    wire [5:0] lut_483_select = {
                             in_data[127],
                             in_data[47],
                             in_data[378],
                             in_data[655],
                             in_data[260],
                             in_data[289]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [63:0] lut_484_table = 64'b0101010001000100010101000100010001010101010101010101010101010101;
    wire [5:0] lut_484_select = {
                             in_data[355],
                             in_data[702],
                             in_data[79],
                             in_data[726],
                             in_data[611],
                             in_data[452]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [63:0] lut_485_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_485_select = {
                             in_data[573],
                             in_data[722],
                             in_data[502],
                             in_data[610],
                             in_data[89],
                             in_data[192]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [63:0] lut_486_table = 64'b1111111100000000111111110010000011111111001000001111111100100010;
    wire [5:0] lut_486_select = {
                             in_data[101],
                             in_data[491],
                             in_data[264],
                             in_data[48],
                             in_data[612],
                             in_data[177]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [63:0] lut_487_table = 64'b0000000011110011000000000111001100000000111100110000000000110011;
    wire [5:0] lut_487_select = {
                             in_data[637],
                             in_data[379],
                             in_data[537],
                             in_data[660],
                             in_data[240],
                             in_data[533]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [63:0] lut_488_table = 64'b0000000000000000000000000000000000000000000000100000000000001111;
    wire [5:0] lut_488_select = {
                             in_data[105],
                             in_data[617],
                             in_data[70],
                             in_data[190],
                             in_data[3],
                             in_data[754]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [63:0] lut_489_table = 64'b1111000000000000111111110100010111110101000001011111110100000101;
    wire [5:0] lut_489_select = {
                             in_data[538],
                             in_data[571],
                             in_data[482],
                             in_data[499],
                             in_data[39],
                             in_data[496]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [63:0] lut_490_table = 64'b1111111111111111111111111111111111111111111111101111111111111110;
    wire [5:0] lut_490_select = {
                             in_data[107],
                             in_data[643],
                             in_data[49],
                             in_data[246],
                             in_data[74],
                             in_data[139]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [63:0] lut_491_table = 64'b1111111111111111000011110000111111111111111111110000111100001100;
    wire [5:0] lut_491_select = {
                             in_data[299],
                             in_data[526],
                             in_data[390],
                             in_data[320],
                             in_data[270],
                             in_data[254]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [63:0] lut_492_table = 64'b0000101100001111001111110000111100000000000000000000001100000000;
    wire [5:0] lut_492_select = {
                             in_data[656],
                             in_data[277],
                             in_data[399],
                             in_data[550],
                             in_data[250],
                             in_data[779]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [63:0] lut_493_table = 64'b0111011101110111011111110111011100000000000000000000000000000000;
    wire [5:0] lut_493_select = {
                             in_data[354],
                             in_data[700],
                             in_data[670],
                             in_data[748],
                             in_data[519],
                             in_data[705]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [63:0] lut_494_table = 64'b0000111111111111000000110000000000001111111111110000001100000000;
    wire [5:0] lut_494_select = {
                             in_data[719],
                             in_data[328],
                             in_data[711],
                             in_data[658],
                             in_data[630],
                             in_data[507]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [63:0] lut_495_table = 64'b0101010111110101010101011111010101000100010101010100010001010101;
    wire [5:0] lut_495_select = {
                             in_data[211],
                             in_data[780],
                             in_data[164],
                             in_data[300],
                             in_data[510],
                             in_data[382]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [63:0] lut_496_table = 64'b0001001100110011001100110011001100000000000100010000000000000001;
    wire [5:0] lut_496_select = {
                             in_data[436],
                             in_data[283],
                             in_data[487],
                             in_data[649],
                             in_data[551],
                             in_data[500]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [63:0] lut_497_table = 64'b0100010000000100010001000000010001010101010101010101010101010101;
    wire [5:0] lut_497_select = {
                             in_data[275],
                             in_data[24],
                             in_data[244],
                             in_data[782],
                             in_data[279],
                             in_data[161]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [63:0] lut_498_table = 64'b0000000000000000000000000000000000000000000000000000001011101111;
    wire [5:0] lut_498_select = {
                             in_data[286],
                             in_data[387],
                             in_data[229],
                             in_data[376],
                             in_data[677],
                             in_data[421]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [63:0] lut_499_table = 64'b1010101010101010111010101111111100101010000000001111101011111111;
    wire [5:0] lut_499_select = {
                             in_data[597],
                             in_data[263],
                             in_data[232],
                             in_data[776],
                             in_data[672],
                             in_data[417]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [63:0] lut_500_table = 64'b1111011111111111000000000000000011111111111101110000000000000000;
    wire [5:0] lut_500_select = {
                             in_data[114],
                             in_data[432],
                             in_data[364],
                             in_data[774],
                             in_data[117],
                             in_data[337]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [63:0] lut_501_table = 64'b0000000000000000000000000000000000000000010101010000000011011111;
    wire [5:0] lut_501_select = {
                             in_data[202],
                             in_data[37],
                             in_data[497],
                             in_data[641],
                             in_data[141],
                             in_data[565]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [63:0] lut_502_table = 64'b1111111111101111010011000100110011111111111011110100110001001100;
    wire [5:0] lut_502_select = {
                             in_data[167],
                             in_data[348],
                             in_data[683],
                             in_data[73],
                             in_data[303],
                             in_data[525]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [63:0] lut_503_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_503_select = {
                             in_data[265],
                             in_data[448],
                             in_data[241],
                             in_data[4],
                             in_data[490],
                             in_data[197]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [63:0] lut_504_table = 64'b1111000011110000111100001111000011111011111100101111101111110010;
    wire [5:0] lut_504_select = {
                             in_data[688],
                             in_data[363],
                             in_data[648],
                             in_data[235],
                             in_data[305],
                             in_data[681]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [63:0] lut_505_table = 64'b0000010100000101000011110000010100000000000000000000000000000000;
    wire [5:0] lut_505_select = {
                             in_data[400],
                             in_data[218],
                             in_data[266],
                             in_data[332],
                             in_data[423],
                             in_data[313]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [63:0] lut_506_table = 64'b1100110011111111000000001100111111001100111111110000000011001111;
    wire [5:0] lut_506_select = {
                             in_data[90],
                             in_data[96],
                             in_data[653],
                             in_data[394],
                             in_data[579],
                             in_data[703]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [63:0] lut_507_table = 64'b1100110011001100111011101110111011101110110011001110111011101110;
    wire [5:0] lut_507_select = {
                             in_data[760],
                             in_data[416],
                             in_data[474],
                             in_data[168],
                             in_data[459],
                             in_data[556]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [63:0] lut_508_table = 64'b1111111111111111111111111111111111101110111011101110111011101110;
    wire [5:0] lut_508_select = {
                             in_data[163],
                             in_data[38],
                             in_data[30],
                             in_data[310],
                             in_data[94],
                             in_data[245]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [63:0] lut_509_table = 64'b1011111100001010101010111010111011111111000010001011101011111110;
    wire [5:0] lut_509_select = {
                             in_data[685],
                             in_data[430],
                             in_data[375],
                             in_data[709],
                             in_data[397],
                             in_data[370]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [63:0] lut_510_table = 64'b1010101000100011101010000010001010001010001100101000100000100010;
    wire [5:0] lut_510_select = {
                             in_data[505],
                             in_data[78],
                             in_data[239],
                             in_data[87],
                             in_data[158],
                             in_data[548]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [63:0] lut_511_table = 64'b1111111111111111111111111111111111111111111111101111111111111110;
    wire [5:0] lut_511_select = {
                             in_data[644],
                             in_data[224],
                             in_data[646],
                             in_data[479],
                             in_data[739],
                             in_data[694]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
    
    // LUT : 512
    wire [63:0] lut_512_table = 64'b1111111111111111111111111111111101010000010100000000000000000000;
    wire [5:0] lut_512_select = {
                             in_data[159],
                             in_data[710],
                             in_data[380],
                             in_data[625],
                             in_data[20],
                             in_data[636]};
    
    wire lut_512_out = lut_512_table[lut_512_select];
    
    generate
    if ( USE_REG ) begin : ff_512
        reg   lut_512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_512_ff <= lut_512_out;
            end
        end
        
        assign out_data[512] = lut_512_ff;
    end
    else begin : no_ff_512
        assign out_data[512] = lut_512_out;
    end
    endgenerate
    
    
    
    // LUT : 513
    wire [63:0] lut_513_table = 64'b0000010100100000101001011010000000000101001000001010011110100000;
    wire [5:0] lut_513_select = {
                             in_data[166],
                             in_data[667],
                             in_data[408],
                             in_data[607],
                             in_data[195],
                             in_data[541]};
    
    wire lut_513_out = lut_513_table[lut_513_select];
    
    generate
    if ( USE_REG ) begin : ff_513
        reg   lut_513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_513_ff <= lut_513_out;
            end
        end
        
        assign out_data[513] = lut_513_ff;
    end
    else begin : no_ff_513
        assign out_data[513] = lut_513_out;
    end
    endgenerate
    
    
    
    // LUT : 514
    wire [63:0] lut_514_table = 64'b1010101000001000111111111010101010101010101010001111111110101010;
    wire [5:0] lut_514_select = {
                             in_data[52],
                             in_data[708],
                             in_data[572],
                             in_data[88],
                             in_data[296],
                             in_data[713]};
    
    wire lut_514_out = lut_514_table[lut_514_select];
    
    generate
    if ( USE_REG ) begin : ff_514
        reg   lut_514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_514_ff <= lut_514_out;
            end
        end
        
        assign out_data[514] = lut_514_ff;
    end
    else begin : no_ff_514
        assign out_data[514] = lut_514_out;
    end
    endgenerate
    
    
    
    // LUT : 515
    wire [63:0] lut_515_table = 64'b0000000000000000000001100000000011101110000000001111111111100111;
    wire [5:0] lut_515_select = {
                             in_data[598],
                             in_data[71],
                             in_data[186],
                             in_data[698],
                             in_data[373],
                             in_data[412]};
    
    wire lut_515_out = lut_515_table[lut_515_select];
    
    generate
    if ( USE_REG ) begin : ff_515
        reg   lut_515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_515_ff <= lut_515_out;
            end
        end
        
        assign out_data[515] = lut_515_ff;
    end
    else begin : no_ff_515
        assign out_data[515] = lut_515_out;
    end
    endgenerate
    
    
    
    // LUT : 516
    wire [63:0] lut_516_table = 64'b0000000000000000000000000000000001010101000000000001000100000000;
    wire [5:0] lut_516_select = {
                             in_data[772],
                             in_data[61],
                             in_data[324],
                             in_data[31],
                             in_data[200],
                             in_data[451]};
    
    wire lut_516_out = lut_516_table[lut_516_select];
    
    generate
    if ( USE_REG ) begin : ff_516
        reg   lut_516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_516_ff <= lut_516_out;
            end
        end
        
        assign out_data[516] = lut_516_ff;
    end
    else begin : no_ff_516
        assign out_data[516] = lut_516_out;
    end
    endgenerate
    
    
    
    // LUT : 517
    wire [63:0] lut_517_table = 64'b1111111110101010111111111110111011111111101010101111111110101010;
    wire [5:0] lut_517_select = {
                             in_data[769],
                             in_data[230],
                             in_data[152],
                             in_data[9],
                             in_data[404],
                             in_data[149]};
    
    wire lut_517_out = lut_517_table[lut_517_select];
    
    generate
    if ( USE_REG ) begin : ff_517
        reg   lut_517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_517_ff <= lut_517_out;
            end
        end
        
        assign out_data[517] = lut_517_ff;
    end
    else begin : no_ff_517
        assign out_data[517] = lut_517_out;
    end
    endgenerate
    
    
    
    // LUT : 518
    wire [63:0] lut_518_table = 64'b1111000011110000001100000011000001111011011111110000000000000000;
    wire [5:0] lut_518_select = {
                             in_data[524],
                             in_data[485],
                             in_data[85],
                             in_data[469],
                             in_data[106],
                             in_data[123]};
    
    wire lut_518_out = lut_518_table[lut_518_select];
    
    generate
    if ( USE_REG ) begin : ff_518
        reg   lut_518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_518_ff <= lut_518_out;
            end
        end
        
        assign out_data[518] = lut_518_ff;
    end
    else begin : no_ff_518
        assign out_data[518] = lut_518_out;
    end
    endgenerate
    
    
    
    // LUT : 519
    wire [63:0] lut_519_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_519_select = {
                             in_data[456],
                             in_data[243],
                             in_data[621],
                             in_data[18],
                             in_data[109],
                             in_data[84]};
    
    wire lut_519_out = lut_519_table[lut_519_select];
    
    generate
    if ( USE_REG ) begin : ff_519
        reg   lut_519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_519_ff <= lut_519_out;
            end
        end
        
        assign out_data[519] = lut_519_ff;
    end
    else begin : no_ff_519
        assign out_data[519] = lut_519_out;
    end
    endgenerate
    
    
    
    // LUT : 520
    wire [63:0] lut_520_table = 64'b1101111101000100111111110100010011111111010101011111111101010101;
    wire [5:0] lut_520_select = {
                             in_data[401],
                             in_data[51],
                             in_data[153],
                             in_data[559],
                             in_data[473],
                             in_data[600]};
    
    wire lut_520_out = lut_520_table[lut_520_select];
    
    generate
    if ( USE_REG ) begin : ff_520
        reg   lut_520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_520_ff <= lut_520_out;
            end
        end
        
        assign out_data[520] = lut_520_ff;
    end
    else begin : no_ff_520
        assign out_data[520] = lut_520_out;
    end
    endgenerate
    
    
    
    // LUT : 521
    wire [63:0] lut_521_table = 64'b1111111111111111111111111111111111111111111111111111111111111100;
    wire [5:0] lut_521_select = {
                             in_data[279],
                             in_data[703],
                             in_data[777],
                             in_data[733],
                             in_data[561],
                             in_data[53]};
    
    wire lut_521_out = lut_521_table[lut_521_select];
    
    generate
    if ( USE_REG ) begin : ff_521
        reg   lut_521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_521_ff <= lut_521_out;
            end
        end
        
        assign out_data[521] = lut_521_ff;
    end
    else begin : no_ff_521
        assign out_data[521] = lut_521_out;
    end
    endgenerate
    
    
    
    // LUT : 522
    wire [63:0] lut_522_table = 64'b0000000000000000000000000000000011110011111100111011001111110011;
    wire [5:0] lut_522_select = {
                             in_data[358],
                             in_data[504],
                             in_data[13],
                             in_data[474],
                             in_data[385],
                             in_data[641]};
    
    wire lut_522_out = lut_522_table[lut_522_select];
    
    generate
    if ( USE_REG ) begin : ff_522
        reg   lut_522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_522_ff <= lut_522_out;
            end
        end
        
        assign out_data[522] = lut_522_ff;
    end
    else begin : no_ff_522
        assign out_data[522] = lut_522_out;
    end
    endgenerate
    
    
    
    // LUT : 523
    wire [63:0] lut_523_table = 64'b1100110011001100110011001100110011011101110011001101110111001100;
    wire [5:0] lut_523_select = {
                             in_data[497],
                             in_data[573],
                             in_data[314],
                             in_data[306],
                             in_data[454],
                             in_data[405]};
    
    wire lut_523_out = lut_523_table[lut_523_select];
    
    generate
    if ( USE_REG ) begin : ff_523
        reg   lut_523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_523_ff <= lut_523_out;
            end
        end
        
        assign out_data[523] = lut_523_ff;
    end
    else begin : no_ff_523
        assign out_data[523] = lut_523_out;
    end
    endgenerate
    
    
    
    // LUT : 524
    wire [63:0] lut_524_table = 64'b1111111111111111101000001010001011111111111111110000000010000000;
    wire [5:0] lut_524_select = {
                             in_data[669],
                             in_data[155],
                             in_data[14],
                             in_data[148],
                             in_data[770],
                             in_data[557]};
    
    wire lut_524_out = lut_524_table[lut_524_select];
    
    generate
    if ( USE_REG ) begin : ff_524
        reg   lut_524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_524_ff <= lut_524_out;
            end
        end
        
        assign out_data[524] = lut_524_ff;
    end
    else begin : no_ff_524
        assign out_data[524] = lut_524_out;
    end
    endgenerate
    
    
    
    // LUT : 525
    wire [63:0] lut_525_table = 64'b0000000000000000000000000000000000001110000001010000111100000101;
    wire [5:0] lut_525_select = {
                             in_data[161],
                             in_data[138],
                             in_data[686],
                             in_data[667],
                             in_data[21],
                             in_data[460]};
    
    wire lut_525_out = lut_525_table[lut_525_select];
    
    generate
    if ( USE_REG ) begin : ff_525
        reg   lut_525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_525_ff <= lut_525_out;
            end
        end
        
        assign out_data[525] = lut_525_ff;
    end
    else begin : no_ff_525
        assign out_data[525] = lut_525_out;
    end
    endgenerate
    
    
    
    // LUT : 526
    wire [63:0] lut_526_table = 64'b0010101100001010101011110000111100101011000000000010111100001000;
    wire [5:0] lut_526_select = {
                             in_data[67],
                             in_data[243],
                             in_data[490],
                             in_data[247],
                             in_data[376],
                             in_data[550]};
    
    wire lut_526_out = lut_526_table[lut_526_select];
    
    generate
    if ( USE_REG ) begin : ff_526
        reg   lut_526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_526_ff <= lut_526_out;
            end
        end
        
        assign out_data[526] = lut_526_ff;
    end
    else begin : no_ff_526
        assign out_data[526] = lut_526_out;
    end
    endgenerate
    
    
    
    // LUT : 527
    wire [63:0] lut_527_table = 64'b0000010100001111000000000000010100000101000011110000000000000111;
    wire [5:0] lut_527_select = {
                             in_data[17],
                             in_data[710],
                             in_data[638],
                             in_data[606],
                             in_data[419],
                             in_data[107]};
    
    wire lut_527_out = lut_527_table[lut_527_select];
    
    generate
    if ( USE_REG ) begin : ff_527
        reg   lut_527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_527_ff <= lut_527_out;
            end
        end
        
        assign out_data[527] = lut_527_ff;
    end
    else begin : no_ff_527
        assign out_data[527] = lut_527_out;
    end
    endgenerate
    
    
    
    // LUT : 528
    wire [63:0] lut_528_table = 64'b1111111111111111111111111111111110111010101110101011101010111010;
    wire [5:0] lut_528_select = {
                             in_data[574],
                             in_data[700],
                             in_data[422],
                             in_data[99],
                             in_data[514],
                             in_data[555]};
    
    wire lut_528_out = lut_528_table[lut_528_select];
    
    generate
    if ( USE_REG ) begin : ff_528
        reg   lut_528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_528_ff <= lut_528_out;
            end
        end
        
        assign out_data[528] = lut_528_ff;
    end
    else begin : no_ff_528
        assign out_data[528] = lut_528_out;
    end
    endgenerate
    
    
    
    // LUT : 529
    wire [63:0] lut_529_table = 64'b1111111111111111111111111111111111111111111110101111111111111010;
    wire [5:0] lut_529_select = {
                             in_data[298],
                             in_data[109],
                             in_data[529],
                             in_data[713],
                             in_data[23],
                             in_data[255]};
    
    wire lut_529_out = lut_529_table[lut_529_select];
    
    generate
    if ( USE_REG ) begin : ff_529
        reg   lut_529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_529_ff <= lut_529_out;
            end
        end
        
        assign out_data[529] = lut_529_ff;
    end
    else begin : no_ff_529
        assign out_data[529] = lut_529_out;
    end
    endgenerate
    
    
    
    // LUT : 530
    wire [63:0] lut_530_table = 64'b1111111111111111111111111111111111111111111111111111111111001100;
    wire [5:0] lut_530_select = {
                             in_data[285],
                             in_data[640],
                             in_data[636],
                             in_data[44],
                             in_data[120],
                             in_data[477]};
    
    wire lut_530_out = lut_530_table[lut_530_select];
    
    generate
    if ( USE_REG ) begin : ff_530
        reg   lut_530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_530_ff <= lut_530_out;
            end
        end
        
        assign out_data[530] = lut_530_ff;
    end
    else begin : no_ff_530
        assign out_data[530] = lut_530_out;
    end
    endgenerate
    
    
    
    // LUT : 531
    wire [63:0] lut_531_table = 64'b1111111111111111111111111111111100000001000001010000000000000001;
    wire [5:0] lut_531_select = {
                             in_data[509],
                             in_data[633],
                             in_data[614],
                             in_data[412],
                             in_data[7],
                             in_data[396]};
    
    wire lut_531_out = lut_531_table[lut_531_select];
    
    generate
    if ( USE_REG ) begin : ff_531
        reg   lut_531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_531_ff <= lut_531_out;
            end
        end
        
        assign out_data[531] = lut_531_ff;
    end
    else begin : no_ff_531
        assign out_data[531] = lut_531_out;
    end
    endgenerate
    
    
    
    // LUT : 532
    wire [63:0] lut_532_table = 64'b0000000000000000111111111111111100000000000000001111111111111111;
    wire [5:0] lut_532_select = {
                             in_data[235],
                             in_data[513],
                             in_data[371],
                             in_data[167],
                             in_data[558],
                             in_data[4]};
    
    wire lut_532_out = lut_532_table[lut_532_select];
    
    generate
    if ( USE_REG ) begin : ff_532
        reg   lut_532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_532_ff <= lut_532_out;
            end
        end
        
        assign out_data[532] = lut_532_ff;
    end
    else begin : no_ff_532
        assign out_data[532] = lut_532_out;
    end
    endgenerate
    
    
    
    // LUT : 533
    wire [63:0] lut_533_table = 64'b0011000011111111000000000011000011110000111111110010000000110000;
    wire [5:0] lut_533_select = {
                             in_data[172],
                             in_data[597],
                             in_data[173],
                             in_data[45],
                             in_data[714],
                             in_data[119]};
    
    wire lut_533_out = lut_533_table[lut_533_select];
    
    generate
    if ( USE_REG ) begin : ff_533
        reg   lut_533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_533_ff <= lut_533_out;
            end
        end
        
        assign out_data[533] = lut_533_ff;
    end
    else begin : no_ff_533
        assign out_data[533] = lut_533_out;
    end
    endgenerate
    
    
    
    // LUT : 534
    wire [63:0] lut_534_table = 64'b0010001100100010001100110010001000100010001000100011001100100010;
    wire [5:0] lut_534_select = {
                             in_data[5],
                             in_data[206],
                             in_data[404],
                             in_data[3],
                             in_data[301],
                             in_data[217]};
    
    wire lut_534_out = lut_534_table[lut_534_select];
    
    generate
    if ( USE_REG ) begin : ff_534
        reg   lut_534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_534_ff <= lut_534_out;
            end
        end
        
        assign out_data[534] = lut_534_ff;
    end
    else begin : no_ff_534
        assign out_data[534] = lut_534_out;
    end
    endgenerate
    
    
    
    // LUT : 535
    wire [63:0] lut_535_table = 64'b1111111111111111000000001111111100000000111111110000000000000000;
    wire [5:0] lut_535_select = {
                             in_data[244],
                             in_data[593],
                             in_data[635],
                             in_data[169],
                             in_data[673],
                             in_data[725]};
    
    wire lut_535_out = lut_535_table[lut_535_select];
    
    generate
    if ( USE_REG ) begin : ff_535
        reg   lut_535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_535_ff <= lut_535_out;
            end
        end
        
        assign out_data[535] = lut_535_ff;
    end
    else begin : no_ff_535
        assign out_data[535] = lut_535_out;
    end
    endgenerate
    
    
    
    // LUT : 536
    wire [63:0] lut_536_table = 64'b1110111111001100111011111100110011101111110011001111111111001110;
    wire [5:0] lut_536_select = {
                             in_data[761],
                             in_data[718],
                             in_data[519],
                             in_data[771],
                             in_data[688],
                             in_data[194]};
    
    wire lut_536_out = lut_536_table[lut_536_select];
    
    generate
    if ( USE_REG ) begin : ff_536
        reg   lut_536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_536_ff <= lut_536_out;
            end
        end
        
        assign out_data[536] = lut_536_ff;
    end
    else begin : no_ff_536
        assign out_data[536] = lut_536_out;
    end
    endgenerate
    
    
    
    // LUT : 537
    wire [63:0] lut_537_table = 64'b1111111101000100111111110100010011111111010001001111111101000110;
    wire [5:0] lut_537_select = {
                             in_data[253],
                             in_data[393],
                             in_data[333],
                             in_data[530],
                             in_data[494],
                             in_data[342]};
    
    wire lut_537_out = lut_537_table[lut_537_select];
    
    generate
    if ( USE_REG ) begin : ff_537
        reg   lut_537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_537_ff <= lut_537_out;
            end
        end
        
        assign out_data[537] = lut_537_ff;
    end
    else begin : no_ff_537
        assign out_data[537] = lut_537_out;
    end
    endgenerate
    
    
    
    // LUT : 538
    wire [63:0] lut_538_table = 64'b0000000000000000111111111111111100001010000010100011111100111111;
    wire [5:0] lut_538_select = {
                             in_data[551],
                             in_data[466],
                             in_data[390],
                             in_data[351],
                             in_data[227],
                             in_data[540]};
    
    wire lut_538_out = lut_538_table[lut_538_select];
    
    generate
    if ( USE_REG ) begin : ff_538
        reg   lut_538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_538_ff <= lut_538_out;
            end
        end
        
        assign out_data[538] = lut_538_ff;
    end
    else begin : no_ff_538
        assign out_data[538] = lut_538_out;
    end
    endgenerate
    
    
    
    // LUT : 539
    wire [63:0] lut_539_table = 64'b1111111111111111000011110000111100001111000010110000000000000000;
    wire [5:0] lut_539_select = {
                             in_data[541],
                             in_data[426],
                             in_data[757],
                             in_data[632],
                             in_data[705],
                             in_data[31]};
    
    wire lut_539_out = lut_539_table[lut_539_select];
    
    generate
    if ( USE_REG ) begin : ff_539
        reg   lut_539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_539_ff <= lut_539_out;
            end
        end
        
        assign out_data[539] = lut_539_ff;
    end
    else begin : no_ff_539
        assign out_data[539] = lut_539_out;
    end
    endgenerate
    
    
    
    // LUT : 540
    wire [63:0] lut_540_table = 64'b1111111111111111111110101111111110101010111111111000000011111010;
    wire [5:0] lut_540_select = {
                             in_data[40],
                             in_data[444],
                             in_data[736],
                             in_data[470],
                             in_data[642],
                             in_data[162]};
    
    wire lut_540_out = lut_540_table[lut_540_select];
    
    generate
    if ( USE_REG ) begin : ff_540
        reg   lut_540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_540_ff <= lut_540_out;
            end
        end
        
        assign out_data[540] = lut_540_ff;
    end
    else begin : no_ff_540
        assign out_data[540] = lut_540_out;
    end
    endgenerate
    
    
    
    // LUT : 541
    wire [63:0] lut_541_table = 64'b1111101011111111111111111111110110110010111111111011000010000000;
    wire [5:0] lut_541_select = {
                             in_data[453],
                             in_data[408],
                             in_data[296],
                             in_data[395],
                             in_data[457],
                             in_data[359]};
    
    wire lut_541_out = lut_541_table[lut_541_select];
    
    generate
    if ( USE_REG ) begin : ff_541
        reg   lut_541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_541_ff <= lut_541_out;
            end
        end
        
        assign out_data[541] = lut_541_ff;
    end
    else begin : no_ff_541
        assign out_data[541] = lut_541_out;
    end
    endgenerate
    
    
    
    // LUT : 542
    wire [63:0] lut_542_table = 64'b0101010101000100110011001101110101010101010001001100110011011101;
    wire [5:0] lut_542_select = {
                             in_data[15],
                             in_data[349],
                             in_data[488],
                             in_data[37],
                             in_data[543],
                             in_data[379]};
    
    wire lut_542_out = lut_542_table[lut_542_select];
    
    generate
    if ( USE_REG ) begin : ff_542
        reg   lut_542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_542_ff <= lut_542_out;
            end
        end
        
        assign out_data[542] = lut_542_ff;
    end
    else begin : no_ff_542
        assign out_data[542] = lut_542_out;
    end
    endgenerate
    
    
    
    // LUT : 543
    wire [63:0] lut_543_table = 64'b1011111110101110101111111010111010101011001010101010101100101010;
    wire [5:0] lut_543_select = {
                             in_data[199],
                             in_data[448],
                             in_data[462],
                             in_data[368],
                             in_data[441],
                             in_data[327]};
    
    wire lut_543_out = lut_543_table[lut_543_select];
    
    generate
    if ( USE_REG ) begin : ff_543
        reg   lut_543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_543_ff <= lut_543_out;
            end
        end
        
        assign out_data[543] = lut_543_ff;
    end
    else begin : no_ff_543
        assign out_data[543] = lut_543_out;
    end
    endgenerate
    
    
    
    // LUT : 544
    wire [63:0] lut_544_table = 64'b0101110101001101010111010101110100001111010011110101110101001101;
    wire [5:0] lut_544_select = {
                             in_data[249],
                             in_data[281],
                             in_data[752],
                             in_data[521],
                             in_data[527],
                             in_data[322]};
    
    wire lut_544_out = lut_544_table[lut_544_select];
    
    generate
    if ( USE_REG ) begin : ff_544
        reg   lut_544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_544_ff <= lut_544_out;
            end
        end
        
        assign out_data[544] = lut_544_ff;
    end
    else begin : no_ff_544
        assign out_data[544] = lut_544_out;
    end
    endgenerate
    
    
    
    // LUT : 545
    wire [63:0] lut_545_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_545_select = {
                             in_data[476],
                             in_data[12],
                             in_data[589],
                             in_data[370],
                             in_data[213],
                             in_data[94]};
    
    wire lut_545_out = lut_545_table[lut_545_select];
    
    generate
    if ( USE_REG ) begin : ff_545
        reg   lut_545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_545_ff <= lut_545_out;
            end
        end
        
        assign out_data[545] = lut_545_ff;
    end
    else begin : no_ff_545
        assign out_data[545] = lut_545_out;
    end
    endgenerate
    
    
    
    // LUT : 546
    wire [63:0] lut_546_table = 64'b1111111111111101111111011101110111001100110011000000000000000000;
    wire [5:0] lut_546_select = {
                             in_data[299],
                             in_data[373],
                             in_data[38],
                             in_data[49],
                             in_data[242],
                             in_data[417]};
    
    wire lut_546_out = lut_546_table[lut_546_select];
    
    generate
    if ( USE_REG ) begin : ff_546
        reg   lut_546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_546_ff <= lut_546_out;
            end
        end
        
        assign out_data[546] = lut_546_ff;
    end
    else begin : no_ff_546
        assign out_data[546] = lut_546_out;
    end
    endgenerate
    
    
    
    // LUT : 547
    wire [63:0] lut_547_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_547_select = {
                             in_data[318],
                             in_data[225],
                             in_data[450],
                             in_data[2],
                             in_data[278],
                             in_data[414]};
    
    wire lut_547_out = lut_547_table[lut_547_select];
    
    generate
    if ( USE_REG ) begin : ff_547
        reg   lut_547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_547_ff <= lut_547_out;
            end
        end
        
        assign out_data[547] = lut_547_ff;
    end
    else begin : no_ff_547
        assign out_data[547] = lut_547_out;
    end
    endgenerate
    
    
    
    // LUT : 548
    wire [63:0] lut_548_table = 64'b0011001100110011001100111111001100110001001100110011001111110011;
    wire [5:0] lut_548_select = {
                             in_data[696],
                             in_data[582],
                             in_data[357],
                             in_data[277],
                             in_data[292],
                             in_data[780]};
    
    wire lut_548_out = lut_548_table[lut_548_select];
    
    generate
    if ( USE_REG ) begin : ff_548
        reg   lut_548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_548_ff <= lut_548_out;
            end
        end
        
        assign out_data[548] = lut_548_ff;
    end
    else begin : no_ff_548
        assign out_data[548] = lut_548_out;
    end
    endgenerate
    
    
    
    // LUT : 549
    wire [63:0] lut_549_table = 64'b0111010111110101101000101011101011110101111101011010101010110010;
    wire [5:0] lut_549_select = {
                             in_data[617],
                             in_data[241],
                             in_data[493],
                             in_data[240],
                             in_data[92],
                             in_data[297]};
    
    wire lut_549_out = lut_549_table[lut_549_select];
    
    generate
    if ( USE_REG ) begin : ff_549
        reg   lut_549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_549_ff <= lut_549_out;
            end
        end
        
        assign out_data[549] = lut_549_ff;
    end
    else begin : no_ff_549
        assign out_data[549] = lut_549_out;
    end
    endgenerate
    
    
    
    // LUT : 550
    wire [63:0] lut_550_table = 64'b1111111111001101111111111111111111001100000001001111111101001101;
    wire [5:0] lut_550_select = {
                             in_data[501],
                             in_data[384],
                             in_data[147],
                             in_data[479],
                             in_data[622],
                             in_data[528]};
    
    wire lut_550_out = lut_550_table[lut_550_select];
    
    generate
    if ( USE_REG ) begin : ff_550
        reg   lut_550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_550_ff <= lut_550_out;
            end
        end
        
        assign out_data[550] = lut_550_ff;
    end
    else begin : no_ff_550
        assign out_data[550] = lut_550_out;
    end
    endgenerate
    
    
    
    // LUT : 551
    wire [63:0] lut_551_table = 64'b1111111111111111111111111111111111111100111111111111000011111100;
    wire [5:0] lut_551_select = {
                             in_data[160],
                             in_data[525],
                             in_data[435],
                             in_data[680],
                             in_data[689],
                             in_data[704]};
    
    wire lut_551_out = lut_551_table[lut_551_select];
    
    generate
    if ( USE_REG ) begin : ff_551
        reg   lut_551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_551_ff <= lut_551_out;
            end
        end
        
        assign out_data[551] = lut_551_ff;
    end
    else begin : no_ff_551
        assign out_data[551] = lut_551_out;
    end
    endgenerate
    
    
    
    // LUT : 552
    wire [63:0] lut_552_table = 64'b0101011101010111000000010000000101011111010111110000000000000001;
    wire [5:0] lut_552_select = {
                             in_data[246],
                             in_data[133],
                             in_data[674],
                             in_data[332],
                             in_data[250],
                             in_data[291]};
    
    wire lut_552_out = lut_552_table[lut_552_select];
    
    generate
    if ( USE_REG ) begin : ff_552
        reg   lut_552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_552_ff <= lut_552_out;
            end
        end
        
        assign out_data[552] = lut_552_ff;
    end
    else begin : no_ff_552
        assign out_data[552] = lut_552_out;
    end
    endgenerate
    
    
    
    // LUT : 553
    wire [63:0] lut_553_table = 64'b0010001000100010001000100010001000100010001000110010001000100010;
    wire [5:0] lut_553_select = {
                             in_data[730],
                             in_data[142],
                             in_data[562],
                             in_data[694],
                             in_data[679],
                             in_data[273]};
    
    wire lut_553_out = lut_553_table[lut_553_select];
    
    generate
    if ( USE_REG ) begin : ff_553
        reg   lut_553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_553_ff <= lut_553_out;
            end
        end
        
        assign out_data[553] = lut_553_ff;
    end
    else begin : no_ff_553
        assign out_data[553] = lut_553_out;
    end
    endgenerate
    
    
    
    // LUT : 554
    wire [63:0] lut_554_table = 64'b1111111111111111111111111111111100000000000000001111111111111100;
    wire [5:0] lut_554_select = {
                             in_data[566],
                             in_data[707],
                             in_data[168],
                             in_data[309],
                             in_data[533],
                             in_data[445]};
    
    wire lut_554_out = lut_554_table[lut_554_select];
    
    generate
    if ( USE_REG ) begin : ff_554
        reg   lut_554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_554_ff <= lut_554_out;
            end
        end
        
        assign out_data[554] = lut_554_ff;
    end
    else begin : no_ff_554
        assign out_data[554] = lut_554_out;
    end
    endgenerate
    
    
    
    // LUT : 555
    wire [63:0] lut_555_table = 64'b1111101111110010111111111111101011111011111100001111111111111010;
    wire [5:0] lut_555_select = {
                             in_data[701],
                             in_data[166],
                             in_data[744],
                             in_data[664],
                             in_data[418],
                             in_data[340]};
    
    wire lut_555_out = lut_555_table[lut_555_select];
    
    generate
    if ( USE_REG ) begin : ff_555
        reg   lut_555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_555_ff <= lut_555_out;
            end
        end
        
        assign out_data[555] = lut_555_ff;
    end
    else begin : no_ff_555
        assign out_data[555] = lut_555_out;
    end
    endgenerate
    
    
    
    // LUT : 556
    wire [63:0] lut_556_table = 64'b1111111111111111111111111111111111111111111111111010101010100000;
    wire [5:0] lut_556_select = {
                             in_data[186],
                             in_data[130],
                             in_data[719],
                             in_data[536],
                             in_data[65],
                             in_data[495]};
    
    wire lut_556_out = lut_556_table[lut_556_select];
    
    generate
    if ( USE_REG ) begin : ff_556
        reg   lut_556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_556_ff <= lut_556_out;
            end
        end
        
        assign out_data[556] = lut_556_ff;
    end
    else begin : no_ff_556
        assign out_data[556] = lut_556_out;
    end
    endgenerate
    
    
    
    // LUT : 557
    wire [63:0] lut_557_table = 64'b1111111111111111111111111111111111111111111011111111111111101110;
    wire [5:0] lut_557_select = {
                             in_data[724],
                             in_data[85],
                             in_data[135],
                             in_data[60],
                             in_data[583],
                             in_data[100]};
    
    wire lut_557_out = lut_557_table[lut_557_select];
    
    generate
    if ( USE_REG ) begin : ff_557
        reg   lut_557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_557_ff <= lut_557_out;
            end
        end
        
        assign out_data[557] = lut_557_ff;
    end
    else begin : no_ff_557
        assign out_data[557] = lut_557_out;
    end
    endgenerate
    
    
    
    // LUT : 558
    wire [63:0] lut_558_table = 64'b1111110010001100111111001000110011111100000011001111110000001100;
    wire [5:0] lut_558_select = {
                             in_data[402],
                             in_data[54],
                             in_data[268],
                             in_data[128],
                             in_data[378],
                             in_data[212]};
    
    wire lut_558_out = lut_558_table[lut_558_select];
    
    generate
    if ( USE_REG ) begin : ff_558
        reg   lut_558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_558_ff <= lut_558_out;
            end
        end
        
        assign out_data[558] = lut_558_ff;
    end
    else begin : no_ff_558
        assign out_data[558] = lut_558_out;
    end
    endgenerate
    
    
    
    // LUT : 559
    wire [63:0] lut_559_table = 64'b1111111111111111101110101111101011111010111111110000100010101010;
    wire [5:0] lut_559_select = {
                             in_data[443],
                             in_data[690],
                             in_data[538],
                             in_data[579],
                             in_data[41],
                             in_data[482]};
    
    wire lut_559_out = lut_559_table[lut_559_select];
    
    generate
    if ( USE_REG ) begin : ff_559
        reg   lut_559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_559_ff <= lut_559_out;
            end
        end
        
        assign out_data[559] = lut_559_ff;
    end
    else begin : no_ff_559
        assign out_data[559] = lut_559_out;
    end
    endgenerate
    
    
    
    // LUT : 560
    wire [63:0] lut_560_table = 64'b1100110001001100110111011101110001000100010001001100110011001100;
    wire [5:0] lut_560_select = {
                             in_data[723],
                             in_data[548],
                             in_data[364],
                             in_data[756],
                             in_data[429],
                             in_data[123]};
    
    wire lut_560_out = lut_560_table[lut_560_select];
    
    generate
    if ( USE_REG ) begin : ff_560
        reg   lut_560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_560_ff <= lut_560_out;
            end
        end
        
        assign out_data[560] = lut_560_ff;
    end
    else begin : no_ff_560
        assign out_data[560] = lut_560_out;
    end
    endgenerate
    
    
    
    // LUT : 561
    wire [63:0] lut_561_table = 64'b1111111111111111111111101111111011111110111111101111100011111000;
    wire [5:0] lut_561_select = {
                             in_data[215],
                             in_data[415],
                             in_data[70],
                             in_data[542],
                             in_data[136],
                             in_data[678]};
    
    wire lut_561_out = lut_561_table[lut_561_select];
    
    generate
    if ( USE_REG ) begin : ff_561
        reg   lut_561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_561_ff <= lut_561_out;
            end
        end
        
        assign out_data[561] = lut_561_ff;
    end
    else begin : no_ff_561
        assign out_data[561] = lut_561_out;
    end
    endgenerate
    
    
    
    // LUT : 562
    wire [63:0] lut_562_table = 64'b1111111111111111001100110011001111111111111111110011001100110011;
    wire [5:0] lut_562_select = {
                             in_data[449],
                             in_data[745],
                             in_data[760],
                             in_data[308],
                             in_data[407],
                             in_data[776]};
    
    wire lut_562_out = lut_562_table[lut_562_select];
    
    generate
    if ( USE_REG ) begin : ff_562
        reg   lut_562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_562_ff <= lut_562_out;
            end
        end
        
        assign out_data[562] = lut_562_ff;
    end
    else begin : no_ff_562
        assign out_data[562] = lut_562_out;
    end
    endgenerate
    
    
    
    // LUT : 563
    wire [63:0] lut_563_table = 64'b1101110111011101100010000000000011111111111111111000110000001000;
    wire [5:0] lut_563_select = {
                             in_data[734],
                             in_data[461],
                             in_data[360],
                             in_data[423],
                             in_data[621],
                             in_data[329]};
    
    wire lut_563_out = lut_563_table[lut_563_select];
    
    generate
    if ( USE_REG ) begin : ff_563
        reg   lut_563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_563_ff <= lut_563_out;
            end
        end
        
        assign out_data[563] = lut_563_ff;
    end
    else begin : no_ff_563
        assign out_data[563] = lut_563_out;
    end
    endgenerate
    
    
    
    // LUT : 564
    wire [63:0] lut_564_table = 64'b1000110010101100101010001010101010101010101110111010101010111010;
    wire [5:0] lut_564_select = {
                             in_data[498],
                             in_data[122],
                             in_data[506],
                             in_data[569],
                             in_data[567],
                             in_data[455]};
    
    wire lut_564_out = lut_564_table[lut_564_select];
    
    generate
    if ( USE_REG ) begin : ff_564
        reg   lut_564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_564_ff <= lut_564_out;
            end
        end
        
        assign out_data[564] = lut_564_ff;
    end
    else begin : no_ff_564
        assign out_data[564] = lut_564_out;
    end
    endgenerate
    
    
    
    // LUT : 565
    wire [63:0] lut_565_table = 64'b1111011111111111111111111111111100000000110011000000000011001100;
    wire [5:0] lut_565_select = {
                             in_data[425],
                             in_data[502],
                             in_data[708],
                             in_data[63],
                             in_data[372],
                             in_data[197]};
    
    wire lut_565_out = lut_565_table[lut_565_select];
    
    generate
    if ( USE_REG ) begin : ff_565
        reg   lut_565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_565_ff <= lut_565_out;
            end
        end
        
        assign out_data[565] = lut_565_ff;
    end
    else begin : no_ff_565
        assign out_data[565] = lut_565_out;
    end
    endgenerate
    
    
    
    // LUT : 566
    wire [63:0] lut_566_table = 64'b1010101000000000111111110000000010101010000000001111111100000000;
    wire [5:0] lut_566_select = {
                             in_data[59],
                             in_data[205],
                             in_data[468],
                             in_data[531],
                             in_data[742],
                             in_data[272]};
    
    wire lut_566_out = lut_566_table[lut_566_select];
    
    generate
    if ( USE_REG ) begin : ff_566
        reg   lut_566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_566_ff <= lut_566_out;
            end
        end
        
        assign out_data[566] = lut_566_ff;
    end
    else begin : no_ff_566
        assign out_data[566] = lut_566_out;
    end
    endgenerate
    
    
    
    // LUT : 567
    wire [63:0] lut_567_table = 64'b1111000011110000111100001111000011110100111100001111010011110000;
    wire [5:0] lut_567_select = {
                             in_data[264],
                             in_data[88],
                             in_data[183],
                             in_data[524],
                             in_data[388],
                             in_data[492]};
    
    wire lut_567_out = lut_567_table[lut_567_select];
    
    generate
    if ( USE_REG ) begin : ff_567
        reg   lut_567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_567_ff <= lut_567_out;
            end
        end
        
        assign out_data[567] = lut_567_ff;
    end
    else begin : no_ff_567
        assign out_data[567] = lut_567_out;
    end
    endgenerate
    
    
    
    // LUT : 568
    wire [63:0] lut_568_table = 64'b0010111100101111000011110000111100001111001011110000111100001111;
    wire [5:0] lut_568_select = {
                             in_data[112],
                             in_data[76],
                             in_data[438],
                             in_data[601],
                             in_data[157],
                             in_data[439]};
    
    wire lut_568_out = lut_568_table[lut_568_select];
    
    generate
    if ( USE_REG ) begin : ff_568
        reg   lut_568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_568_ff <= lut_568_out;
            end
        end
        
        assign out_data[568] = lut_568_ff;
    end
    else begin : no_ff_568
        assign out_data[568] = lut_568_out;
    end
    endgenerate
    
    
    
    // LUT : 569
    wire [63:0] lut_569_table = 64'b0000000000000000000000010000000100000001000000010010011100100111;
    wire [5:0] lut_569_select = {
                             in_data[326],
                             in_data[229],
                             in_data[749],
                             in_data[545],
                             in_data[339],
                             in_data[259]};
    
    wire lut_569_out = lut_569_table[lut_569_select];
    
    generate
    if ( USE_REG ) begin : ff_569
        reg   lut_569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_569_ff <= lut_569_out;
            end
        end
        
        assign out_data[569] = lut_569_ff;
    end
    else begin : no_ff_569
        assign out_data[569] = lut_569_out;
    end
    endgenerate
    
    
    
    // LUT : 570
    wire [63:0] lut_570_table = 64'b1111111100001010111111110000000011111111100010101111111100000000;
    wire [5:0] lut_570_select = {
                             in_data[9],
                             in_data[68],
                             in_data[374],
                             in_data[475],
                             in_data[113],
                             in_data[275]};
    
    wire lut_570_out = lut_570_table[lut_570_select];
    
    generate
    if ( USE_REG ) begin : ff_570
        reg   lut_570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_570_ff <= lut_570_out;
            end
        end
        
        assign out_data[570] = lut_570_ff;
    end
    else begin : no_ff_570
        assign out_data[570] = lut_570_out;
    end
    endgenerate
    
    
    
    // LUT : 571
    wire [63:0] lut_571_table = 64'b0101110101010101010101010101010101000100010001000100010001000100;
    wire [5:0] lut_571_select = {
                             in_data[300],
                             in_data[591],
                             in_data[544],
                             in_data[767],
                             in_data[687],
                             in_data[434]};
    
    wire lut_571_out = lut_571_table[lut_571_select];
    
    generate
    if ( USE_REG ) begin : ff_571
        reg   lut_571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_571_ff <= lut_571_out;
            end
        end
        
        assign out_data[571] = lut_571_ff;
    end
    else begin : no_ff_571
        assign out_data[571] = lut_571_out;
    end
    endgenerate
    
    
    
    // LUT : 572
    wire [63:0] lut_572_table = 64'b0001000000000000000000000000000001010101010101010101010001010000;
    wire [5:0] lut_572_select = {
                             in_data[537],
                             in_data[549],
                             in_data[615],
                             in_data[338],
                             in_data[295],
                             in_data[684]};
    
    wire lut_572_out = lut_572_table[lut_572_select];
    
    generate
    if ( USE_REG ) begin : ff_572
        reg   lut_572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_572_ff <= lut_572_out;
            end
        end
        
        assign out_data[572] = lut_572_ff;
    end
    else begin : no_ff_572
        assign out_data[572] = lut_572_out;
    end
    endgenerate
    
    
    
    // LUT : 573
    wire [63:0] lut_573_table = 64'b1111111111111111111111111111111111111101100011001111110100000000;
    wire [5:0] lut_573_select = {
                             in_data[575],
                             in_data[198],
                             in_data[584],
                             in_data[383],
                             in_data[552],
                             in_data[702]};
    
    wire lut_573_out = lut_573_table[lut_573_select];
    
    generate
    if ( USE_REG ) begin : ff_573
        reg   lut_573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_573_ff <= lut_573_out;
            end
        end
        
        assign out_data[573] = lut_573_ff;
    end
    else begin : no_ff_573
        assign out_data[573] = lut_573_out;
    end
    endgenerate
    
    
    
    // LUT : 574
    wire [63:0] lut_574_table = 64'b1011001011110000101100101111000000001010111100000000101011110000;
    wire [5:0] lut_574_select = {
                             in_data[293],
                             in_data[84],
                             in_data[177],
                             in_data[483],
                             in_data[263],
                             in_data[345]};
    
    wire lut_574_out = lut_574_table[lut_574_select];
    
    generate
    if ( USE_REG ) begin : ff_574
        reg   lut_574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_574_ff <= lut_574_out;
            end
        end
        
        assign out_data[574] = lut_574_ff;
    end
    else begin : no_ff_574
        assign out_data[574] = lut_574_out;
    end
    endgenerate
    
    
    
    // LUT : 575
    wire [63:0] lut_575_table = 64'b0000001100110011001000110011001100010011001100110001001100110011;
    wire [5:0] lut_575_select = {
                             in_data[252],
                             in_data[18],
                             in_data[467],
                             in_data[739],
                             in_data[324],
                             in_data[740]};
    
    wire lut_575_out = lut_575_table[lut_575_select];
    
    generate
    if ( USE_REG ) begin : ff_575
        reg   lut_575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_575_ff <= lut_575_out;
            end
        end
        
        assign out_data[575] = lut_575_ff;
    end
    else begin : no_ff_575
        assign out_data[575] = lut_575_out;
    end
    endgenerate
    
    
    
    // LUT : 576
    wire [63:0] lut_576_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_576_select = {
                             in_data[489],
                             in_data[754],
                             in_data[728],
                             in_data[682],
                             in_data[697],
                             in_data[81]};
    
    wire lut_576_out = lut_576_table[lut_576_select];
    
    generate
    if ( USE_REG ) begin : ff_576
        reg   lut_576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_576_ff <= lut_576_out;
            end
        end
        
        assign out_data[576] = lut_576_ff;
    end
    else begin : no_ff_576
        assign out_data[576] = lut_576_out;
    end
    endgenerate
    
    
    
    // LUT : 577
    wire [63:0] lut_577_table = 64'b1011111110101010111111111111101011111111000010101111111110101111;
    wire [5:0] lut_577_select = {
                             in_data[353],
                             in_data[102],
                             in_data[218],
                             in_data[628],
                             in_data[392],
                             in_data[623]};
    
    wire lut_577_out = lut_577_table[lut_577_select];
    
    generate
    if ( USE_REG ) begin : ff_577
        reg   lut_577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_577_ff <= lut_577_out;
            end
        end
        
        assign out_data[577] = lut_577_ff;
    end
    else begin : no_ff_577
        assign out_data[577] = lut_577_out;
    end
    endgenerate
    
    
    
    // LUT : 578
    wire [63:0] lut_578_table = 64'b1111111000001000111111100000100011111111100011101111111110001110;
    wire [5:0] lut_578_select = {
                             in_data[311],
                             in_data[22],
                             in_data[608],
                             in_data[656],
                             in_data[485],
                             in_data[305]};
    
    wire lut_578_out = lut_578_table[lut_578_select];
    
    generate
    if ( USE_REG ) begin : ff_578
        reg   lut_578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_578_ff <= lut_578_out;
            end
        end
        
        assign out_data[578] = lut_578_ff;
    end
    else begin : no_ff_578
        assign out_data[578] = lut_578_out;
    end
    endgenerate
    
    
    
    // LUT : 579
    wire [63:0] lut_579_table = 64'b0000000011010101000000000100000011101010111111111111111111111111;
    wire [5:0] lut_579_select = {
                             in_data[465],
                             in_data[224],
                             in_data[346],
                             in_data[699],
                             in_data[95],
                             in_data[207]};
    
    wire lut_579_out = lut_579_table[lut_579_select];
    
    generate
    if ( USE_REG ) begin : ff_579
        reg   lut_579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_579_ff <= lut_579_out;
            end
        end
        
        assign out_data[579] = lut_579_ff;
    end
    else begin : no_ff_579
        assign out_data[579] = lut_579_out;
    end
    endgenerate
    
    
    
    // LUT : 580
    wire [63:0] lut_580_table = 64'b0011101110111011101110111011101111111111111111111010101110101010;
    wire [5:0] lut_580_select = {
                             in_data[625],
                             in_data[565],
                             in_data[334],
                             in_data[440],
                             in_data[380],
                             in_data[96]};
    
    wire lut_580_out = lut_580_table[lut_580_select];
    
    generate
    if ( USE_REG ) begin : ff_580
        reg   lut_580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_580_ff <= lut_580_out;
            end
        end
        
        assign out_data[580] = lut_580_ff;
    end
    else begin : no_ff_580
        assign out_data[580] = lut_580_out;
    end
    endgenerate
    
    
    
    // LUT : 581
    wire [63:0] lut_581_table = 64'b1111111111111111111111111111111111101010111010101110101011111010;
    wire [5:0] lut_581_select = {
                             in_data[151],
                             in_data[580],
                             in_data[27],
                             in_data[683],
                             in_data[262],
                             in_data[121]};
    
    wire lut_581_out = lut_581_table[lut_581_select];
    
    generate
    if ( USE_REG ) begin : ff_581
        reg   lut_581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_581_ff <= lut_581_out;
            end
        end
        
        assign out_data[581] = lut_581_ff;
    end
    else begin : no_ff_581
        assign out_data[581] = lut_581_out;
    end
    endgenerate
    
    
    
    // LUT : 582
    wire [63:0] lut_582_table = 64'b0000010100000101000001010000010100000101000001010000010100000101;
    wire [5:0] lut_582_select = {
                             in_data[643],
                             in_data[768],
                             in_data[775],
                             in_data[261],
                             in_data[646],
                             in_data[594]};
    
    wire lut_582_out = lut_582_table[lut_582_select];
    
    generate
    if ( USE_REG ) begin : ff_582
        reg   lut_582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_582_ff <= lut_582_out;
            end
        end
        
        assign out_data[582] = lut_582_ff;
    end
    else begin : no_ff_582
        assign out_data[582] = lut_582_out;
    end
    endgenerate
    
    
    
    // LUT : 583
    wire [63:0] lut_583_table = 64'b1111111111111111001010100010101011111111111111110010101000001010;
    wire [5:0] lut_583_select = {
                             in_data[751],
                             in_data[491],
                             in_data[79],
                             in_data[534],
                             in_data[698],
                             in_data[663]};
    
    wire lut_583_out = lut_583_table[lut_583_select];
    
    generate
    if ( USE_REG ) begin : ff_583
        reg   lut_583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_583_ff <= lut_583_out;
            end
        end
        
        assign out_data[583] = lut_583_ff;
    end
    else begin : no_ff_583
        assign out_data[583] = lut_583_out;
    end
    endgenerate
    
    
    
    // LUT : 584
    wire [63:0] lut_584_table = 64'b0000000000000000000000000000000010101010101010101111111111111111;
    wire [5:0] lut_584_select = {
                             in_data[269],
                             in_data[657],
                             in_data[39],
                             in_data[766],
                             in_data[114],
                             in_data[712]};
    
    wire lut_584_out = lut_584_table[lut_584_select];
    
    generate
    if ( USE_REG ) begin : ff_584
        reg   lut_584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_584_ff <= lut_584_out;
            end
        end
        
        assign out_data[584] = lut_584_ff;
    end
    else begin : no_ff_584
        assign out_data[584] = lut_584_out;
    end
    endgenerate
    
    
    
    // LUT : 585
    wire [63:0] lut_585_table = 64'b1111111110101111111011111010111111111111001011111111111100111111;
    wire [5:0] lut_585_select = {
                             in_data[189],
                             in_data[753],
                             in_data[499],
                             in_data[209],
                             in_data[381],
                             in_data[362]};
    
    wire lut_585_out = lut_585_table[lut_585_select];
    
    generate
    if ( USE_REG ) begin : ff_585
        reg   lut_585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_585_ff <= lut_585_out;
            end
        end
        
        assign out_data[585] = lut_585_ff;
    end
    else begin : no_ff_585
        assign out_data[585] = lut_585_out;
    end
    endgenerate
    
    
    
    // LUT : 586
    wire [63:0] lut_586_table = 64'b1100100011001000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_586_select = {
                             in_data[350],
                             in_data[176],
                             in_data[336],
                             in_data[738],
                             in_data[331],
                             in_data[458]};
    
    wire lut_586_out = lut_586_table[lut_586_select];
    
    generate
    if ( USE_REG ) begin : ff_586
        reg   lut_586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_586_ff <= lut_586_out;
            end
        end
        
        assign out_data[586] = lut_586_ff;
    end
    else begin : no_ff_586
        assign out_data[586] = lut_586_out;
    end
    endgenerate
    
    
    
    // LUT : 587
    wire [63:0] lut_587_table = 64'b0000000000000000101000101010000001010101000101001111111111111111;
    wire [5:0] lut_587_select = {
                             in_data[188],
                             in_data[321],
                             in_data[764],
                             in_data[203],
                             in_data[639],
                             in_data[546]};
    
    wire lut_587_out = lut_587_table[lut_587_select];
    
    generate
    if ( USE_REG ) begin : ff_587
        reg   lut_587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_587_ff <= lut_587_out;
            end
        end
        
        assign out_data[587] = lut_587_ff;
    end
    else begin : no_ff_587
        assign out_data[587] = lut_587_out;
    end
    endgenerate
    
    
    
    // LUT : 588
    wire [63:0] lut_588_table = 64'b0000000000000000000000000000000001000000010100001111000011110010;
    wire [5:0] lut_588_select = {
                             in_data[662],
                             in_data[146],
                             in_data[62],
                             in_data[317],
                             in_data[722],
                             in_data[230]};
    
    wire lut_588_out = lut_588_table[lut_588_select];
    
    generate
    if ( USE_REG ) begin : ff_588
        reg   lut_588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_588_ff <= lut_588_out;
            end
        end
        
        assign out_data[588] = lut_588_ff;
    end
    else begin : no_ff_588
        assign out_data[588] = lut_588_out;
    end
    endgenerate
    
    
    
    // LUT : 589
    wire [63:0] lut_589_table = 64'b0000000000000000000000000000000011111111111111001111111111110000;
    wire [5:0] lut_589_select = {
                             in_data[741],
                             in_data[563],
                             in_data[73],
                             in_data[400],
                             in_data[46],
                             in_data[50]};
    
    wire lut_589_out = lut_589_table[lut_589_select];
    
    generate
    if ( USE_REG ) begin : ff_589
        reg   lut_589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_589_ff <= lut_589_out;
            end
        end
        
        assign out_data[589] = lut_589_ff;
    end
    else begin : no_ff_589
        assign out_data[589] = lut_589_out;
    end
    endgenerate
    
    
    
    // LUT : 590
    wire [63:0] lut_590_table = 64'b1111111111111111101110110000001111001100010101010010001000000000;
    wire [5:0] lut_590_select = {
                             in_data[179],
                             in_data[572],
                             in_data[553],
                             in_data[772],
                             in_data[510],
                             in_data[211]};
    
    wire lut_590_out = lut_590_table[lut_590_select];
    
    generate
    if ( USE_REG ) begin : ff_590
        reg   lut_590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_590_ff <= lut_590_out;
            end
        end
        
        assign out_data[590] = lut_590_ff;
    end
    else begin : no_ff_590
        assign out_data[590] = lut_590_out;
    end
    endgenerate
    
    
    
    // LUT : 591
    wire [63:0] lut_591_table = 64'b0000000000000000000000000000000000000000111111110000000011111111;
    wire [5:0] lut_591_select = {
                             in_data[377],
                             in_data[196],
                             in_data[182],
                             in_data[118],
                             in_data[143],
                             in_data[420]};
    
    wire lut_591_out = lut_591_table[lut_591_select];
    
    generate
    if ( USE_REG ) begin : ff_591
        reg   lut_591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_591_ff <= lut_591_out;
            end
        end
        
        assign out_data[591] = lut_591_ff;
    end
    else begin : no_ff_591
        assign out_data[591] = lut_591_out;
    end
    endgenerate
    
    
    
    // LUT : 592
    wire [63:0] lut_592_table = 64'b0010101010101010000010101010101000101010101010100010101010101111;
    wire [5:0] lut_592_select = {
                             in_data[695],
                             in_data[214],
                             in_data[451],
                             in_data[556],
                             in_data[586],
                             in_data[220]};
    
    wire lut_592_out = lut_592_table[lut_592_select];
    
    generate
    if ( USE_REG ) begin : ff_592
        reg   lut_592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_592_ff <= lut_592_out;
            end
        end
        
        assign out_data[592] = lut_592_ff;
    end
    else begin : no_ff_592
        assign out_data[592] = lut_592_out;
    end
    endgenerate
    
    
    
    // LUT : 593
    wire [63:0] lut_593_table = 64'b0000001100000011001111110000101100000000000000000000000000000000;
    wire [5:0] lut_593_select = {
                             in_data[433],
                             in_data[303],
                             in_data[672],
                             in_data[629],
                             in_data[190],
                             in_data[590]};
    
    wire lut_593_out = lut_593_table[lut_593_select];
    
    generate
    if ( USE_REG ) begin : ff_593
        reg   lut_593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_593_ff <= lut_593_out;
            end
        end
        
        assign out_data[593] = lut_593_ff;
    end
    else begin : no_ff_593
        assign out_data[593] = lut_593_out;
    end
    endgenerate
    
    
    
    // LUT : 594
    wire [63:0] lut_594_table = 64'b0001000100010001001101110011011100010000000100010011001100010011;
    wire [5:0] lut_594_select = {
                             in_data[221],
                             in_data[399],
                             in_data[782],
                             in_data[313],
                             in_data[398],
                             in_data[204]};
    
    wire lut_594_out = lut_594_table[lut_594_select];
    
    generate
    if ( USE_REG ) begin : ff_594
        reg   lut_594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_594_ff <= lut_594_out;
            end
        end
        
        assign out_data[594] = lut_594_ff;
    end
    else begin : no_ff_594
        assign out_data[594] = lut_594_out;
    end
    endgenerate
    
    
    
    // LUT : 595
    wire [63:0] lut_595_table = 64'b0000000000000000011101110110000000000000000000001111111101110001;
    wire [5:0] lut_595_select = {
                             in_data[709],
                             in_data[348],
                             in_data[236],
                             in_data[11],
                             in_data[496],
                             in_data[294]};
    
    wire lut_595_out = lut_595_table[lut_595_select];
    
    generate
    if ( USE_REG ) begin : ff_595
        reg   lut_595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_595_ff <= lut_595_out;
            end
        end
        
        assign out_data[595] = lut_595_ff;
    end
    else begin : no_ff_595
        assign out_data[595] = lut_595_out;
    end
    endgenerate
    
    
    
    // LUT : 596
    wire [63:0] lut_596_table = 64'b0000000000000000111111111111111100000000000000001111111111111111;
    wire [5:0] lut_596_select = {
                             in_data[32],
                             in_data[347],
                             in_data[30],
                             in_data[644],
                             in_data[517],
                             in_data[778]};
    
    wire lut_596_out = lut_596_table[lut_596_select];
    
    generate
    if ( USE_REG ) begin : ff_596
        reg   lut_596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_596_ff <= lut_596_out;
            end
        end
        
        assign out_data[596] = lut_596_ff;
    end
    else begin : no_ff_596
        assign out_data[596] = lut_596_out;
    end
    endgenerate
    
    
    
    // LUT : 597
    wire [63:0] lut_597_table = 64'b1000110011001110100011001000110011001100110011101100110010001100;
    wire [5:0] lut_597_select = {
                             in_data[337],
                             in_data[452],
                             in_data[316],
                             in_data[387],
                             in_data[430],
                             in_data[578]};
    
    wire lut_597_out = lut_597_table[lut_597_select];
    
    generate
    if ( USE_REG ) begin : ff_597
        reg   lut_597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_597_ff <= lut_597_out;
            end
        end
        
        assign out_data[597] = lut_597_ff;
    end
    else begin : no_ff_597
        assign out_data[597] = lut_597_out;
    end
    endgenerate
    
    
    
    // LUT : 598
    wire [63:0] lut_598_table = 64'b0011001111110000001100110111000000100010111111100010001011111111;
    wire [5:0] lut_598_select = {
                             in_data[436],
                             in_data[36],
                             in_data[302],
                             in_data[369],
                             in_data[596],
                             in_data[127]};
    
    wire lut_598_out = lut_598_table[lut_598_select];
    
    generate
    if ( USE_REG ) begin : ff_598
        reg   lut_598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_598_ff <= lut_598_out;
            end
        end
        
        assign out_data[598] = lut_598_ff;
    end
    else begin : no_ff_598
        assign out_data[598] = lut_598_out;
    end
    endgenerate
    
    
    
    // LUT : 599
    wire [63:0] lut_599_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_599_select = {
                             in_data[150],
                             in_data[200],
                             in_data[487],
                             in_data[671],
                             in_data[187],
                             in_data[238]};
    
    wire lut_599_out = lut_599_table[lut_599_select];
    
    generate
    if ( USE_REG ) begin : ff_599
        reg   lut_599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_599_ff <= lut_599_out;
            end
        end
        
        assign out_data[599] = lut_599_ff;
    end
    else begin : no_ff_599
        assign out_data[599] = lut_599_out;
    end
    endgenerate
    
    
    
    // LUT : 600
    wire [63:0] lut_600_table = 64'b0101010101010101010101110101011100000000000000000000000000000000;
    wire [5:0] lut_600_select = {
                             in_data[343],
                             in_data[386],
                             in_data[232],
                             in_data[620],
                             in_data[354],
                             in_data[652]};
    
    wire lut_600_out = lut_600_table[lut_600_select];
    
    generate
    if ( USE_REG ) begin : ff_600
        reg   lut_600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_600_ff <= lut_600_out;
            end
        end
        
        assign out_data[600] = lut_600_ff;
    end
    else begin : no_ff_600
        assign out_data[600] = lut_600_out;
    end
    endgenerate
    
    
    
    // LUT : 601
    wire [63:0] lut_601_table = 64'b1010111010101010111011101010101011101110111011101111111011101110;
    wire [5:0] lut_601_select = {
                             in_data[774],
                             in_data[505],
                             in_data[676],
                             in_data[781],
                             in_data[320],
                             in_data[653]};
    
    wire lut_601_out = lut_601_table[lut_601_select];
    
    generate
    if ( USE_REG ) begin : ff_601
        reg   lut_601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_601_ff <= lut_601_out;
            end
        end
        
        assign out_data[601] = lut_601_ff;
    end
    else begin : no_ff_601
        assign out_data[601] = lut_601_out;
    end
    endgenerate
    
    
    
    // LUT : 602
    wire [63:0] lut_602_table = 64'b0000000000000000000000000000000010101010101010101010101010101010;
    wire [5:0] lut_602_select = {
                             in_data[271],
                             in_data[731],
                             in_data[222],
                             in_data[180],
                             in_data[692],
                             in_data[516]};
    
    wire lut_602_out = lut_602_table[lut_602_select];
    
    generate
    if ( USE_REG ) begin : ff_602
        reg   lut_602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_602_ff <= lut_602_out;
            end
        end
        
        assign out_data[602] = lut_602_ff;
    end
    else begin : no_ff_602
        assign out_data[602] = lut_602_out;
    end
    endgenerate
    
    
    
    // LUT : 603
    wire [63:0] lut_603_table = 64'b1111111111111111111111111111111101010101111111111100110011111110;
    wire [5:0] lut_603_select = {
                             in_data[715],
                             in_data[603],
                             in_data[598],
                             in_data[64],
                             in_data[675],
                             in_data[237]};
    
    wire lut_603_out = lut_603_table[lut_603_select];
    
    generate
    if ( USE_REG ) begin : ff_603
        reg   lut_603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_603_ff <= lut_603_out;
            end
        end
        
        assign out_data[603] = lut_603_ff;
    end
    else begin : no_ff_603
        assign out_data[603] = lut_603_out;
    end
    endgenerate
    
    
    
    // LUT : 604
    wire [63:0] lut_604_table = 64'b0011001100110011001100110111001100110011001100110011001100110011;
    wire [5:0] lut_604_select = {
                             in_data[685],
                             in_data[735],
                             in_data[406],
                             in_data[69],
                             in_data[270],
                             in_data[91]};
    
    wire lut_604_out = lut_604_table[lut_604_select];
    
    generate
    if ( USE_REG ) begin : ff_604
        reg   lut_604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_604_ff <= lut_604_out;
            end
        end
        
        assign out_data[604] = lut_604_ff;
    end
    else begin : no_ff_604
        assign out_data[604] = lut_604_out;
    end
    endgenerate
    
    
    
    // LUT : 605
    wire [63:0] lut_605_table = 64'b0101011100010101010101010000010101010111000101010101011100000001;
    wire [5:0] lut_605_select = {
                             in_data[57],
                             in_data[446],
                             in_data[693],
                             in_data[71],
                             in_data[595],
                             in_data[156]};
    
    wire lut_605_out = lut_605_table[lut_605_select];
    
    generate
    if ( USE_REG ) begin : ff_605
        reg   lut_605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_605_ff <= lut_605_out;
            end
        end
        
        assign out_data[605] = lut_605_ff;
    end
    else begin : no_ff_605
        assign out_data[605] = lut_605_out;
    end
    endgenerate
    
    
    
    // LUT : 606
    wire [63:0] lut_606_table = 64'b1111111111111111111011111010111100001111001011110000010000000101;
    wire [5:0] lut_606_select = {
                             in_data[658],
                             in_data[284],
                             in_data[58],
                             in_data[612],
                             in_data[755],
                             in_data[459]};
    
    wire lut_606_out = lut_606_table[lut_606_select];
    
    generate
    if ( USE_REG ) begin : ff_606
        reg   lut_606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_606_ff <= lut_606_out;
            end
        end
        
        assign out_data[606] = lut_606_ff;
    end
    else begin : no_ff_606
        assign out_data[606] = lut_606_out;
    end
    endgenerate
    
    
    
    // LUT : 607
    wire [63:0] lut_607_table = 64'b1111111111111111111111111111111111111100111011001111110011101100;
    wire [5:0] lut_607_select = {
                             in_data[634],
                             in_data[115],
                             in_data[428],
                             in_data[154],
                             in_data[260],
                             in_data[66]};
    
    wire lut_607_out = lut_607_table[lut_607_select];
    
    generate
    if ( USE_REG ) begin : ff_607
        reg   lut_607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_607_ff <= lut_607_out;
            end
        end
        
        assign out_data[607] = lut_607_ff;
    end
    else begin : no_ff_607
        assign out_data[607] = lut_607_out;
    end
    endgenerate
    
    
    
    // LUT : 608
    wire [63:0] lut_608_table = 64'b1010101010101010101010101010101010101111101011101010111110101111;
    wire [5:0] lut_608_select = {
                             in_data[464],
                             in_data[56],
                             in_data[108],
                             in_data[231],
                             in_data[52],
                             in_data[126]};
    
    wire lut_608_out = lut_608_table[lut_608_select];
    
    generate
    if ( USE_REG ) begin : ff_608
        reg   lut_608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_608_ff <= lut_608_out;
            end
        end
        
        assign out_data[608] = lut_608_ff;
    end
    else begin : no_ff_608
        assign out_data[608] = lut_608_out;
    end
    endgenerate
    
    
    
    // LUT : 609
    wire [63:0] lut_609_table = 64'b1111111111111111111111111111111111111111111111101111111111111110;
    wire [5:0] lut_609_select = {
                             in_data[330],
                             in_data[410],
                             in_data[257],
                             in_data[43],
                             in_data[747],
                             in_data[310]};
    
    wire lut_609_out = lut_609_table[lut_609_select];
    
    generate
    if ( USE_REG ) begin : ff_609
        reg   lut_609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_609_ff <= lut_609_out;
            end
        end
        
        assign out_data[609] = lut_609_ff;
    end
    else begin : no_ff_609
        assign out_data[609] = lut_609_out;
    end
    endgenerate
    
    
    
    // LUT : 610
    wire [63:0] lut_610_table = 64'b0000000010000000000000000000000010001111111011110000111100000111;
    wire [5:0] lut_610_select = {
                             in_data[152],
                             in_data[500],
                             in_data[547],
                             in_data[508],
                             in_data[605],
                             in_data[604]};
    
    wire lut_610_out = lut_610_table[lut_610_select];
    
    generate
    if ( USE_REG ) begin : ff_610
        reg   lut_610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_610_ff <= lut_610_out;
            end
        end
        
        assign out_data[610] = lut_610_ff;
    end
    else begin : no_ff_610
        assign out_data[610] = lut_610_out;
    end
    endgenerate
    
    
    
    // LUT : 611
    wire [63:0] lut_611_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_611_select = {
                             in_data[363],
                             in_data[391],
                             in_data[323],
                             in_data[290],
                             in_data[280],
                             in_data[145]};
    
    wire lut_611_out = lut_611_table[lut_611_select];
    
    generate
    if ( USE_REG ) begin : ff_611
        reg   lut_611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_611_ff <= lut_611_out;
            end
        end
        
        assign out_data[611] = lut_611_ff;
    end
    else begin : no_ff_611
        assign out_data[611] = lut_611_out;
    end
    endgenerate
    
    
    
    // LUT : 612
    wire [63:0] lut_612_table = 64'b0000111101011111000010101010101000001111010111110000101010101010;
    wire [5:0] lut_612_select = {
                             in_data[48],
                             in_data[581],
                             in_data[184],
                             in_data[131],
                             in_data[140],
                             in_data[512]};
    
    wire lut_612_out = lut_612_table[lut_612_select];
    
    generate
    if ( USE_REG ) begin : ff_612
        reg   lut_612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_612_ff <= lut_612_out;
            end
        end
        
        assign out_data[612] = lut_612_ff;
    end
    else begin : no_ff_612
        assign out_data[612] = lut_612_out;
    end
    endgenerate
    
    
    
    // LUT : 613
    wire [63:0] lut_613_table = 64'b1010101010101010000000000010001010101010101010101000000010101010;
    wire [5:0] lut_613_select = {
                             in_data[424],
                             in_data[219],
                             in_data[607],
                             in_data[616],
                             in_data[750],
                             in_data[515]};
    
    wire lut_613_out = lut_613_table[lut_613_select];
    
    generate
    if ( USE_REG ) begin : ff_613
        reg   lut_613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_613_ff <= lut_613_out;
            end
        end
        
        assign out_data[613] = lut_613_ff;
    end
    else begin : no_ff_613
        assign out_data[613] = lut_613_out;
    end
    endgenerate
    
    
    
    // LUT : 614
    wire [63:0] lut_614_table = 64'b1111111101110101111111111111110101010101010101000101010101010101;
    wire [5:0] lut_614_select = {
                             in_data[248],
                             in_data[783],
                             in_data[307],
                             in_data[627],
                             in_data[25],
                             in_data[382]};
    
    wire lut_614_out = lut_614_table[lut_614_select];
    
    generate
    if ( USE_REG ) begin : ff_614
        reg   lut_614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_614_ff <= lut_614_out;
            end
        end
        
        assign out_data[614] = lut_614_ff;
    end
    else begin : no_ff_614
        assign out_data[614] = lut_614_out;
    end
    endgenerate
    
    
    
    // LUT : 615
    wire [63:0] lut_615_table = 64'b0011000000000000000100000000000011110011000010111111001100001111;
    wire [5:0] lut_615_select = {
                             in_data[403],
                             in_data[765],
                             in_data[522],
                             in_data[375],
                             in_data[312],
                             in_data[82]};
    
    wire lut_615_out = lut_615_table[lut_615_select];
    
    generate
    if ( USE_REG ) begin : ff_615
        reg   lut_615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_615_ff <= lut_615_out;
            end
        end
        
        assign out_data[615] = lut_615_ff;
    end
    else begin : no_ff_615
        assign out_data[615] = lut_615_out;
    end
    endgenerate
    
    
    
    // LUT : 616
    wire [63:0] lut_616_table = 64'b1111111111111111111111111111000011111111111111111111101111110000;
    wire [5:0] lut_616_select = {
                             in_data[437],
                             in_data[288],
                             in_data[163],
                             in_data[341],
                             in_data[758],
                             in_data[727]};
    
    wire lut_616_out = lut_616_table[lut_616_select];
    
    generate
    if ( USE_REG ) begin : ff_616
        reg   lut_616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_616_ff <= lut_616_out;
            end
        end
        
        assign out_data[616] = lut_616_ff;
    end
    else begin : no_ff_616
        assign out_data[616] = lut_616_out;
    end
    endgenerate
    
    
    
    // LUT : 617
    wire [63:0] lut_617_table = 64'b0000000011111111000000001111111100000000111101010000000011110101;
    wire [5:0] lut_617_select = {
                             in_data[471],
                             in_data[34],
                             in_data[159],
                             in_data[0],
                             in_data[647],
                             in_data[746]};
    
    wire lut_617_out = lut_617_table[lut_617_select];
    
    generate
    if ( USE_REG ) begin : ff_617
        reg   lut_617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_617_ff <= lut_617_out;
            end
        end
        
        assign out_data[617] = lut_617_ff;
    end
    else begin : no_ff_617
        assign out_data[617] = lut_617_out;
    end
    endgenerate
    
    
    
    // LUT : 618
    wire [63:0] lut_618_table = 64'b0010101000101010001010100010101000101011001010110010101100101011;
    wire [5:0] lut_618_select = {
                             in_data[599],
                             in_data[335],
                             in_data[16],
                             in_data[175],
                             in_data[134],
                             in_data[304]};
    
    wire lut_618_out = lut_618_table[lut_618_select];
    
    generate
    if ( USE_REG ) begin : ff_618
        reg   lut_618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_618_ff <= lut_618_out;
            end
        end
        
        assign out_data[618] = lut_618_ff;
    end
    else begin : no_ff_618
        assign out_data[618] = lut_618_out;
    end
    endgenerate
    
    
    
    // LUT : 619
    wire [63:0] lut_619_table = 64'b1100110011001100110011111100111111001100110011001100111111001111;
    wire [5:0] lut_619_select = {
                             in_data[26],
                             in_data[149],
                             in_data[421],
                             in_data[315],
                             in_data[681],
                             in_data[732]};
    
    wire lut_619_out = lut_619_table[lut_619_select];
    
    generate
    if ( USE_REG ) begin : ff_619
        reg   lut_619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_619_ff <= lut_619_out;
            end
        end
        
        assign out_data[619] = lut_619_ff;
    end
    else begin : no_ff_619
        assign out_data[619] = lut_619_out;
    end
    endgenerate
    
    
    
    // LUT : 620
    wire [63:0] lut_620_table = 64'b0001000100010001000100010001000100010001000100010001000100010001;
    wire [5:0] lut_620_select = {
                             in_data[98],
                             in_data[144],
                             in_data[762],
                             in_data[78],
                             in_data[356],
                             in_data[716]};
    
    wire lut_620_out = lut_620_table[lut_620_select];
    
    generate
    if ( USE_REG ) begin : ff_620
        reg   lut_620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_620_ff <= lut_620_out;
            end
        end
        
        assign out_data[620] = lut_620_ff;
    end
    else begin : no_ff_620
        assign out_data[620] = lut_620_out;
    end
    endgenerate
    
    
    
    // LUT : 621
    wire [63:0] lut_621_table = 64'b0100010111010101000000000000010011010101110101010000010100000101;
    wire [5:0] lut_621_select = {
                             in_data[367],
                             in_data[361],
                             in_data[394],
                             in_data[463],
                             in_data[192],
                             in_data[245]};
    
    wire lut_621_out = lut_621_table[lut_621_select];
    
    generate
    if ( USE_REG ) begin : ff_621
        reg   lut_621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_621_ff <= lut_621_out;
            end
        end
        
        assign out_data[621] = lut_621_ff;
    end
    else begin : no_ff_621
        assign out_data[621] = lut_621_out;
    end
    endgenerate
    
    
    
    // LUT : 622
    wire [63:0] lut_622_table = 64'b0000000000000000000000000001000100000000101010100000000001110111;
    wire [5:0] lut_622_select = {
                             in_data[106],
                             in_data[654],
                             in_data[185],
                             in_data[223],
                             in_data[254],
                             in_data[568]};
    
    wire lut_622_out = lut_622_table[lut_622_select];
    
    generate
    if ( USE_REG ) begin : ff_622
        reg   lut_622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_622_ff <= lut_622_out;
            end
        end
        
        assign out_data[622] = lut_622_ff;
    end
    else begin : no_ff_622
        assign out_data[622] = lut_622_out;
    end
    endgenerate
    
    
    
    // LUT : 623
    wire [63:0] lut_623_table = 64'b1111111111111111111111111010101011111111111111111111111110101010;
    wire [5:0] lut_623_select = {
                             in_data[47],
                             in_data[178],
                             in_data[389],
                             in_data[626],
                             in_data[6],
                             in_data[472]};
    
    wire lut_623_out = lut_623_table[lut_623_select];
    
    generate
    if ( USE_REG ) begin : ff_623
        reg   lut_623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_623_ff <= lut_623_out;
            end
        end
        
        assign out_data[623] = lut_623_ff;
    end
    else begin : no_ff_623
        assign out_data[623] = lut_623_out;
    end
    endgenerate
    
    
    
    // LUT : 624
    wire [63:0] lut_624_table = 64'b1111111111111111101010101011101011111111111111111010101010101010;
    wire [5:0] lut_624_select = {
                             in_data[28],
                             in_data[743],
                             in_data[587],
                             in_data[560],
                             in_data[283],
                             in_data[287]};
    
    wire lut_624_out = lut_624_table[lut_624_select];
    
    generate
    if ( USE_REG ) begin : ff_624
        reg   lut_624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_624_ff <= lut_624_out;
            end
        end
        
        assign out_data[624] = lut_624_ff;
    end
    else begin : no_ff_624
        assign out_data[624] = lut_624_out;
    end
    endgenerate
    
    
    
    // LUT : 625
    wire [63:0] lut_625_table = 64'b0111000101110001011100010111000101110001011100010101000101110001;
    wire [5:0] lut_625_select = {
                             in_data[86],
                             in_data[588],
                             in_data[773],
                             in_data[691],
                             in_data[210],
                             in_data[539]};
    
    wire lut_625_out = lut_625_table[lut_625_select];
    
    generate
    if ( USE_REG ) begin : ff_625
        reg   lut_625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_625_ff <= lut_625_out;
            end
        end
        
        assign out_data[625] = lut_625_ff;
    end
    else begin : no_ff_625
        assign out_data[625] = lut_625_out;
    end
    endgenerate
    
    
    
    // LUT : 626
    wire [63:0] lut_626_table = 64'b1111111111111010111111111010101011111111111110101111111110101010;
    wire [5:0] lut_626_select = {
                             in_data[42],
                             in_data[366],
                             in_data[325],
                             in_data[585],
                             in_data[666],
                             in_data[650]};
    
    wire lut_626_out = lut_626_table[lut_626_select];
    
    generate
    if ( USE_REG ) begin : ff_626
        reg   lut_626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_626_ff <= lut_626_out;
            end
        end
        
        assign out_data[626] = lut_626_ff;
    end
    else begin : no_ff_626
        assign out_data[626] = lut_626_out;
    end
    endgenerate
    
    
    
    // LUT : 627
    wire [63:0] lut_627_table = 64'b1111111111111111111111111111111111111111101110101111111110101010;
    wire [5:0] lut_627_select = {
                             in_data[105],
                             in_data[170],
                             in_data[174],
                             in_data[645],
                             in_data[729],
                             in_data[648]};
    
    wire lut_627_out = lut_627_table[lut_627_select];
    
    generate
    if ( USE_REG ) begin : ff_627
        reg   lut_627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_627_ff <= lut_627_out;
            end
        end
        
        assign out_data[627] = lut_627_ff;
    end
    else begin : no_ff_627
        assign out_data[627] = lut_627_out;
    end
    endgenerate
    
    
    
    // LUT : 628
    wire [63:0] lut_628_table = 64'b0000000011111111000000001111111100100000111111110000000011111111;
    wire [5:0] lut_628_select = {
                             in_data[216],
                             in_data[75],
                             in_data[442],
                             in_data[611],
                             in_data[90],
                             in_data[258]};
    
    wire lut_628_out = lut_628_table[lut_628_select];
    
    generate
    if ( USE_REG ) begin : ff_628
        reg   lut_628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_628_ff <= lut_628_out;
            end
        end
        
        assign out_data[628] = lut_628_ff;
    end
    else begin : no_ff_628
        assign out_data[628] = lut_628_out;
    end
    endgenerate
    
    
    
    // LUT : 629
    wire [63:0] lut_629_table = 64'b1111111111001100111111111101110011111111110011001111111111001100;
    wire [5:0] lut_629_select = {
                             in_data[478],
                             in_data[365],
                             in_data[132],
                             in_data[89],
                             in_data[413],
                             in_data[523]};
    
    wire lut_629_out = lut_629_table[lut_629_select];
    
    generate
    if ( USE_REG ) begin : ff_629
        reg   lut_629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_629_ff <= lut_629_out;
            end
        end
        
        assign out_data[629] = lut_629_ff;
    end
    else begin : no_ff_629
        assign out_data[629] = lut_629_out;
    end
    endgenerate
    
    
    
    // LUT : 630
    wire [63:0] lut_630_table = 64'b0000000000000000010101010101010100000000000000000101010101010101;
    wire [5:0] lut_630_select = {
                             in_data[195],
                             in_data[193],
                             in_data[116],
                             in_data[267],
                             in_data[171],
                             in_data[520]};
    
    wire lut_630_out = lut_630_table[lut_630_select];
    
    generate
    if ( USE_REG ) begin : ff_630
        reg   lut_630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_630_ff <= lut_630_out;
            end
        end
        
        assign out_data[630] = lut_630_ff;
    end
    else begin : no_ff_630
        assign out_data[630] = lut_630_out;
    end
    endgenerate
    
    
    
    // LUT : 631
    wire [63:0] lut_631_table = 64'b1011101111111111101110111011101100010001000000000001000100000000;
    wire [5:0] lut_631_select = {
                             in_data[234],
                             in_data[637],
                             in_data[651],
                             in_data[226],
                             in_data[481],
                             in_data[631]};
    
    wire lut_631_out = lut_631_table[lut_631_select];
    
    generate
    if ( USE_REG ) begin : ff_631
        reg   lut_631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_631_ff <= lut_631_out;
            end
        end
        
        assign out_data[631] = lut_631_ff;
    end
    else begin : no_ff_631
        assign out_data[631] = lut_631_out;
    end
    endgenerate
    
    
    
    // LUT : 632
    wire [63:0] lut_632_table = 64'b1111111111111111111111011111110111110100111111111111010011111101;
    wire [5:0] lut_632_select = {
                             in_data[748],
                             in_data[609],
                             in_data[411],
                             in_data[711],
                             in_data[706],
                             in_data[137]};
    
    wire lut_632_out = lut_632_table[lut_632_select];
    
    generate
    if ( USE_REG ) begin : ff_632
        reg   lut_632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_632_ff <= lut_632_out;
            end
        end
        
        assign out_data[632] = lut_632_ff;
    end
    else begin : no_ff_632
        assign out_data[632] = lut_632_out;
    end
    endgenerate
    
    
    
    // LUT : 633
    wire [63:0] lut_633_table = 64'b1010101010101010101010101010101010101010101011111010101010101111;
    wire [5:0] lut_633_select = {
                             in_data[77],
                             in_data[33],
                             in_data[484],
                             in_data[649],
                             in_data[613],
                             in_data[129]};
    
    wire lut_633_out = lut_633_table[lut_633_select];
    
    generate
    if ( USE_REG ) begin : ff_633
        reg   lut_633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_633_ff <= lut_633_out;
            end
        end
        
        assign out_data[633] = lut_633_ff;
    end
    else begin : no_ff_633
        assign out_data[633] = lut_633_out;
    end
    endgenerate
    
    
    
    // LUT : 634
    wire [63:0] lut_634_table = 64'b1111111110101111101010100000000011111111111111111111111110101010;
    wire [5:0] lut_634_select = {
                             in_data[164],
                             in_data[660],
                             in_data[432],
                             in_data[201],
                             in_data[111],
                             in_data[526]};
    
    wire lut_634_out = lut_634_table[lut_634_select];
    
    generate
    if ( USE_REG ) begin : ff_634
        reg   lut_634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_634_ff <= lut_634_out;
            end
        end
        
        assign out_data[634] = lut_634_ff;
    end
    else begin : no_ff_634
        assign out_data[634] = lut_634_out;
    end
    endgenerate
    
    
    
    // LUT : 635
    wire [63:0] lut_635_table = 64'b1010101010101010111111101111111110101010101010101111111111111111;
    wire [5:0] lut_635_select = {
                             in_data[665],
                             in_data[266],
                             in_data[165],
                             in_data[191],
                             in_data[117],
                             in_data[125]};
    
    wire lut_635_out = lut_635_table[lut_635_select];
    
    generate
    if ( USE_REG ) begin : ff_635
        reg   lut_635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_635_ff <= lut_635_out;
            end
        end
        
        assign out_data[635] = lut_635_ff;
    end
    else begin : no_ff_635
        assign out_data[635] = lut_635_out;
    end
    endgenerate
    
    
    
    // LUT : 636
    wire [63:0] lut_636_table = 64'b0011000000110011000100000011001100000000001100110000000000110001;
    wire [5:0] lut_636_select = {
                             in_data[35],
                             in_data[276],
                             in_data[677],
                             in_data[564],
                             in_data[737],
                             in_data[1]};
    
    wire lut_636_out = lut_636_table[lut_636_select];
    
    generate
    if ( USE_REG ) begin : ff_636
        reg   lut_636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_636_ff <= lut_636_out;
            end
        end
        
        assign out_data[636] = lut_636_ff;
    end
    else begin : no_ff_636
        assign out_data[636] = lut_636_out;
    end
    endgenerate
    
    
    
    // LUT : 637
    wire [63:0] lut_637_table = 64'b0101000000000001010101010101010101010000000001010111010101010101;
    wire [5:0] lut_637_select = {
                             in_data[110],
                             in_data[456],
                             in_data[624],
                             in_data[239],
                             in_data[10],
                             in_data[469]};
    
    wire lut_637_out = lut_637_table[lut_637_select];
    
    generate
    if ( USE_REG ) begin : ff_637
        reg   lut_637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_637_ff <= lut_637_out;
            end
        end
        
        assign out_data[637] = lut_637_ff;
    end
    else begin : no_ff_637
        assign out_data[637] = lut_637_out;
    end
    endgenerate
    
    
    
    // LUT : 638
    wire [63:0] lut_638_table = 64'b0000000000000100000000000000010000000000000000110000000000000011;
    wire [5:0] lut_638_select = {
                             in_data[431],
                             in_data[87],
                             in_data[202],
                             in_data[717],
                             in_data[409],
                             in_data[72]};
    
    wire lut_638_out = lut_638_table[lut_638_select];
    
    generate
    if ( USE_REG ) begin : ff_638
        reg   lut_638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_638_ff <= lut_638_out;
            end
        end
        
        assign out_data[638] = lut_638_ff;
    end
    else begin : no_ff_638
        assign out_data[638] = lut_638_out;
    end
    endgenerate
    
    
    
    // LUT : 639
    wire [63:0] lut_639_table = 64'b1111000111110001011100000101000011110001111100010101000001010000;
    wire [5:0] lut_639_select = {
                             in_data[779],
                             in_data[721],
                             in_data[8],
                             in_data[427],
                             in_data[282],
                             in_data[256]};
    
    wire lut_639_out = lut_639_table[lut_639_select];
    
    generate
    if ( USE_REG ) begin : ff_639
        reg   lut_639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_639_ff <= lut_639_out;
            end
        end
        
        assign out_data[639] = lut_639_ff;
    end
    else begin : no_ff_639
        assign out_data[639] = lut_639_out;
    end
    endgenerate
    
    
    
    // LUT : 640
    wire [63:0] lut_640_table = 64'b0000000000000000000000000000000000001011000011110000001100000011;
    wire [5:0] lut_640_select = {
                             in_data[720],
                             in_data[618],
                             in_data[61],
                             in_data[103],
                             in_data[352],
                             in_data[251]};
    
    wire lut_640_out = lut_640_table[lut_640_select];
    
    generate
    if ( USE_REG ) begin : ff_640
        reg   lut_640_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_640_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_640_ff <= lut_640_out;
            end
        end
        
        assign out_data[640] = lut_640_ff;
    end
    else begin : no_ff_640
        assign out_data[640] = lut_640_out;
    end
    endgenerate
    
    
    
    // LUT : 641
    wire [63:0] lut_641_table = 64'b1111111111011001111111010101000011111111110111011111110111010000;
    wire [5:0] lut_641_select = {
                             in_data[726],
                             in_data[93],
                             in_data[511],
                             in_data[554],
                             in_data[181],
                             in_data[158]};
    
    wire lut_641_out = lut_641_table[lut_641_select];
    
    generate
    if ( USE_REG ) begin : ff_641
        reg   lut_641_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_641_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_641_ff <= lut_641_out;
            end
        end
        
        assign out_data[641] = lut_641_ff;
    end
    else begin : no_ff_641
        assign out_data[641] = lut_641_out;
    end
    endgenerate
    
    
    
    // LUT : 642
    wire [63:0] lut_642_table = 64'b1111010001110100111100000011000011111110011111111111110000111111;
    wire [5:0] lut_642_select = {
                             in_data[659],
                             in_data[480],
                             in_data[486],
                             in_data[576],
                             in_data[630],
                             in_data[319]};
    
    wire lut_642_out = lut_642_table[lut_642_select];
    
    generate
    if ( USE_REG ) begin : ff_642
        reg   lut_642_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_642_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_642_ff <= lut_642_out;
            end
        end
        
        assign out_data[642] = lut_642_ff;
    end
    else begin : no_ff_642
        assign out_data[642] = lut_642_out;
    end
    endgenerate
    
    
    
    // LUT : 643
    wire [63:0] lut_643_table = 64'b1111111111101110111111111110111011111111111011101111111111101110;
    wire [5:0] lut_643_select = {
                             in_data[507],
                             in_data[532],
                             in_data[228],
                             in_data[55],
                             in_data[124],
                             in_data[655]};
    
    wire lut_643_out = lut_643_table[lut_643_select];
    
    generate
    if ( USE_REG ) begin : ff_643
        reg   lut_643_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_643_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_643_ff <= lut_643_out;
            end
        end
        
        assign out_data[643] = lut_643_ff;
    end
    else begin : no_ff_643
        assign out_data[643] = lut_643_out;
    end
    endgenerate
    
    
    
    // LUT : 644
    wire [63:0] lut_644_table = 64'b1111000001110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_644_select = {
                             in_data[619],
                             in_data[104],
                             in_data[759],
                             in_data[328],
                             in_data[74],
                             in_data[289]};
    
    wire lut_644_out = lut_644_table[lut_644_select];
    
    generate
    if ( USE_REG ) begin : ff_644
        reg   lut_644_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_644_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_644_ff <= lut_644_out;
            end
        end
        
        assign out_data[644] = lut_644_ff;
    end
    else begin : no_ff_644
        assign out_data[644] = lut_644_out;
    end
    endgenerate
    
    
    
    // LUT : 645
    wire [63:0] lut_645_table = 64'b0101111111011111010101010101010101011111010111110000010101010101;
    wire [5:0] lut_645_select = {
                             in_data[97],
                             in_data[274],
                             in_data[535],
                             in_data[602],
                             in_data[80],
                             in_data[208]};
    
    wire lut_645_out = lut_645_table[lut_645_select];
    
    generate
    if ( USE_REG ) begin : ff_645
        reg   lut_645_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_645_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_645_ff <= lut_645_out;
            end
        end
        
        assign out_data[645] = lut_645_ff;
    end
    else begin : no_ff_645
        assign out_data[645] = lut_645_out;
    end
    endgenerate
    
    
    
    // LUT : 646
    wire [63:0] lut_646_table = 64'b1111000011110000111110001111100011110000111100001111110011111100;
    wire [5:0] lut_646_select = {
                             in_data[83],
                             in_data[518],
                             in_data[503],
                             in_data[344],
                             in_data[101],
                             in_data[24]};
    
    wire lut_646_out = lut_646_table[lut_646_select];
    
    generate
    if ( USE_REG ) begin : ff_646
        reg   lut_646_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_646_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_646_ff <= lut_646_out;
            end
        end
        
        assign out_data[646] = lut_646_ff;
    end
    else begin : no_ff_646
        assign out_data[646] = lut_646_out;
    end
    endgenerate
    
    
    
    // LUT : 647
    wire [63:0] lut_647_table = 64'b0000000000000000000000000101010100000000000000000000000001010101;
    wire [5:0] lut_647_select = {
                             in_data[763],
                             in_data[416],
                             in_data[661],
                             in_data[139],
                             in_data[141],
                             in_data[610]};
    
    wire lut_647_out = lut_647_table[lut_647_select];
    
    generate
    if ( USE_REG ) begin : ff_647
        reg   lut_647_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_647_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_647_ff <= lut_647_out;
            end
        end
        
        assign out_data[647] = lut_647_ff;
    end
    else begin : no_ff_647
        assign out_data[647] = lut_647_out;
    end
    endgenerate
    
    
    
    // LUT : 648
    wire [63:0] lut_648_table = 64'b0000000000100010001000100010001100000000001110110000000000110011;
    wire [5:0] lut_648_select = {
                             in_data[570],
                             in_data[286],
                             in_data[571],
                             in_data[447],
                             in_data[592],
                             in_data[668]};
    
    wire lut_648_out = lut_648_table[lut_648_select];
    
    generate
    if ( USE_REG ) begin : ff_648
        reg   lut_648_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_648_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_648_ff <= lut_648_out;
            end
        end
        
        assign out_data[648] = lut_648_ff;
    end
    else begin : no_ff_648
        assign out_data[648] = lut_648_out;
    end
    endgenerate
    
    
    
    // LUT : 649
    wire [63:0] lut_649_table = 64'b0000000100000101000010100000011100001111000011110010111100001111;
    wire [5:0] lut_649_select = {
                             in_data[233],
                             in_data[355],
                             in_data[29],
                             in_data[577],
                             in_data[769],
                             in_data[397]};
    
    wire lut_649_out = lut_649_table[lut_649_select];
    
    generate
    if ( USE_REG ) begin : ff_649
        reg   lut_649_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_649_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_649_ff <= lut_649_out;
            end
        end
        
        assign out_data[649] = lut_649_ff;
    end
    else begin : no_ff_649
        assign out_data[649] = lut_649_out;
    end
    endgenerate
    
    
    
    // LUT : 650
    wire [63:0] lut_650_table = 64'b0000000000000000000010111010111100000000000000001111111111111111;
    wire [5:0] lut_650_select = {
                             in_data[232],
                             in_data[518],
                             in_data[20],
                             in_data[670],
                             in_data[265],
                             in_data[19]};
    
    wire lut_650_out = lut_650_table[lut_650_select];
    
    generate
    if ( USE_REG ) begin : ff_650
        reg   lut_650_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_650_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_650_ff <= lut_650_out;
            end
        end
        
        assign out_data[650] = lut_650_ff;
    end
    else begin : no_ff_650
        assign out_data[650] = lut_650_out;
    end
    endgenerate
    
    
    
    // LUT : 651
    wire [63:0] lut_651_table = 64'b1101110111111101110111001101110011111101111111011101110011001100;
    wire [5:0] lut_651_select = {
                             in_data[695],
                             in_data[625],
                             in_data[634],
                             in_data[709],
                             in_data[267],
                             in_data[597]};
    
    wire lut_651_out = lut_651_table[lut_651_select];
    
    generate
    if ( USE_REG ) begin : ff_651
        reg   lut_651_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_651_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_651_ff <= lut_651_out;
            end
        end
        
        assign out_data[651] = lut_651_ff;
    end
    else begin : no_ff_651
        assign out_data[651] = lut_651_out;
    end
    endgenerate
    
    
    
    // LUT : 652
    wire [63:0] lut_652_table = 64'b1111110011111100111111001111111011000000111111001100000011111100;
    wire [5:0] lut_652_select = {
                             in_data[495],
                             in_data[641],
                             in_data[575],
                             in_data[456],
                             in_data[494],
                             in_data[42]};
    
    wire lut_652_out = lut_652_table[lut_652_select];
    
    generate
    if ( USE_REG ) begin : ff_652
        reg   lut_652_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_652_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_652_ff <= lut_652_out;
            end
        end
        
        assign out_data[652] = lut_652_ff;
    end
    else begin : no_ff_652
        assign out_data[652] = lut_652_out;
    end
    endgenerate
    
    
    
    // LUT : 653
    wire [63:0] lut_653_table = 64'b1101110111001100110011001100110011011101010011001100110011001100;
    wire [5:0] lut_653_select = {
                             in_data[770],
                             in_data[154],
                             in_data[524],
                             in_data[4],
                             in_data[437],
                             in_data[256]};
    
    wire lut_653_out = lut_653_table[lut_653_select];
    
    generate
    if ( USE_REG ) begin : ff_653
        reg   lut_653_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_653_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_653_ff <= lut_653_out;
            end
        end
        
        assign out_data[653] = lut_653_ff;
    end
    else begin : no_ff_653
        assign out_data[653] = lut_653_out;
    end
    endgenerate
    
    
    
    // LUT : 654
    wire [63:0] lut_654_table = 64'b1011111100000000111111110000000010101010101110111010101010111011;
    wire [5:0] lut_654_select = {
                             in_data[512],
                             in_data[647],
                             in_data[301],
                             in_data[731],
                             in_data[204],
                             in_data[608]};
    
    wire lut_654_out = lut_654_table[lut_654_select];
    
    generate
    if ( USE_REG ) begin : ff_654
        reg   lut_654_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_654_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_654_ff <= lut_654_out;
            end
        end
        
        assign out_data[654] = lut_654_ff;
    end
    else begin : no_ff_654
        assign out_data[654] = lut_654_out;
    end
    endgenerate
    
    
    
    // LUT : 655
    wire [63:0] lut_655_table = 64'b0111011100000000011100110000000001110011000000000111001100000000;
    wire [5:0] lut_655_select = {
                             in_data[773],
                             in_data[728],
                             in_data[213],
                             in_data[183],
                             in_data[149],
                             in_data[122]};
    
    wire lut_655_out = lut_655_table[lut_655_select];
    
    generate
    if ( USE_REG ) begin : ff_655
        reg   lut_655_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_655_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_655_ff <= lut_655_out;
            end
        end
        
        assign out_data[655] = lut_655_ff;
    end
    else begin : no_ff_655
        assign out_data[655] = lut_655_out;
    end
    endgenerate
    
    
    
    // LUT : 656
    wire [63:0] lut_656_table = 64'b0000010100000101010001010000010101010101000001010000010100000000;
    wire [5:0] lut_656_select = {
                             in_data[384],
                             in_data[548],
                             in_data[352],
                             in_data[94],
                             in_data[422],
                             in_data[545]};
    
    wire lut_656_out = lut_656_table[lut_656_select];
    
    generate
    if ( USE_REG ) begin : ff_656
        reg   lut_656_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_656_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_656_ff <= lut_656_out;
            end
        end
        
        assign out_data[656] = lut_656_ff;
    end
    else begin : no_ff_656
        assign out_data[656] = lut_656_out;
    end
    endgenerate
    
    
    
    // LUT : 657
    wire [63:0] lut_657_table = 64'b1111111111110011000000111010001011111111111110111010101110110011;
    wire [5:0] lut_657_select = {
                             in_data[145],
                             in_data[473],
                             in_data[315],
                             in_data[292],
                             in_data[656],
                             in_data[637]};
    
    wire lut_657_out = lut_657_table[lut_657_select];
    
    generate
    if ( USE_REG ) begin : ff_657
        reg   lut_657_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_657_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_657_ff <= lut_657_out;
            end
        end
        
        assign out_data[657] = lut_657_ff;
    end
    else begin : no_ff_657
        assign out_data[657] = lut_657_out;
    end
    endgenerate
    
    
    
    // LUT : 658
    wire [63:0] lut_658_table = 64'b0000000011111111010000001111111100000000000000000000000000000101;
    wire [5:0] lut_658_select = {
                             in_data[513],
                             in_data[452],
                             in_data[326],
                             in_data[50],
                             in_data[110],
                             in_data[13]};
    
    wire lut_658_out = lut_658_table[lut_658_select];
    
    generate
    if ( USE_REG ) begin : ff_658
        reg   lut_658_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_658_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_658_ff <= lut_658_out;
            end
        end
        
        assign out_data[658] = lut_658_ff;
    end
    else begin : no_ff_658
        assign out_data[658] = lut_658_out;
    end
    endgenerate
    
    
    
    // LUT : 659
    wire [63:0] lut_659_table = 64'b1111111111001111111111111111111111001111110011111100111111001111;
    wire [5:0] lut_659_select = {
                             in_data[203],
                             in_data[115],
                             in_data[138],
                             in_data[603],
                             in_data[133],
                             in_data[393]};
    
    wire lut_659_out = lut_659_table[lut_659_select];
    
    generate
    if ( USE_REG ) begin : ff_659
        reg   lut_659_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_659_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_659_ff <= lut_659_out;
            end
        end
        
        assign out_data[659] = lut_659_ff;
    end
    else begin : no_ff_659
        assign out_data[659] = lut_659_out;
    end
    endgenerate
    
    
    
    // LUT : 660
    wire [63:0] lut_660_table = 64'b1111110011111100111111001111110011101100111011001111110011111100;
    wire [5:0] lut_660_select = {
                             in_data[611],
                             in_data[275],
                             in_data[17],
                             in_data[537],
                             in_data[485],
                             in_data[638]};
    
    wire lut_660_out = lut_660_table[lut_660_select];
    
    generate
    if ( USE_REG ) begin : ff_660
        reg   lut_660_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_660_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_660_ff <= lut_660_out;
            end
        end
        
        assign out_data[660] = lut_660_ff;
    end
    else begin : no_ff_660
        assign out_data[660] = lut_660_out;
    end
    endgenerate
    
    
    
    // LUT : 661
    wire [63:0] lut_661_table = 64'b0001000100010001000100010001000100010001000100010001000100010001;
    wire [5:0] lut_661_select = {
                             in_data[8],
                             in_data[226],
                             in_data[617],
                             in_data[642],
                             in_data[233],
                             in_data[380]};
    
    wire lut_661_out = lut_661_table[lut_661_select];
    
    generate
    if ( USE_REG ) begin : ff_661
        reg   lut_661_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_661_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_661_ff <= lut_661_out;
            end
        end
        
        assign out_data[661] = lut_661_ff;
    end
    else begin : no_ff_661
        assign out_data[661] = lut_661_out;
    end
    endgenerate
    
    
    
    // LUT : 662
    wire [63:0] lut_662_table = 64'b1101110111111111110011001100110011011101111111011100110011101100;
    wire [5:0] lut_662_select = {
                             in_data[58],
                             in_data[211],
                             in_data[108],
                             in_data[766],
                             in_data[706],
                             in_data[102]};
    
    wire lut_662_out = lut_662_table[lut_662_select];
    
    generate
    if ( USE_REG ) begin : ff_662
        reg   lut_662_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_662_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_662_ff <= lut_662_out;
            end
        end
        
        assign out_data[662] = lut_662_ff;
    end
    else begin : no_ff_662
        assign out_data[662] = lut_662_out;
    end
    endgenerate
    
    
    
    // LUT : 663
    wire [63:0] lut_663_table = 64'b1111111111111111111111111101111100000000000000000000110100001101;
    wire [5:0] lut_663_select = {
                             in_data[397],
                             in_data[509],
                             in_data[755],
                             in_data[97],
                             in_data[475],
                             in_data[46]};
    
    wire lut_663_out = lut_663_table[lut_663_select];
    
    generate
    if ( USE_REG ) begin : ff_663
        reg   lut_663_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_663_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_663_ff <= lut_663_out;
            end
        end
        
        assign out_data[663] = lut_663_ff;
    end
    else begin : no_ff_663
        assign out_data[663] = lut_663_out;
    end
    endgenerate
    
    
    
    // LUT : 664
    wire [63:0] lut_664_table = 64'b0010001000100010101010101010101011111111111111111110111011111110;
    wire [5:0] lut_664_select = {
                             in_data[543],
                             in_data[493],
                             in_data[26],
                             in_data[36],
                             in_data[436],
                             in_data[746]};
    
    wire lut_664_out = lut_664_table[lut_664_select];
    
    generate
    if ( USE_REG ) begin : ff_664
        reg   lut_664_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_664_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_664_ff <= lut_664_out;
            end
        end
        
        assign out_data[664] = lut_664_ff;
    end
    else begin : no_ff_664
        assign out_data[664] = lut_664_out;
    end
    endgenerate
    
    
    
    // LUT : 665
    wire [63:0] lut_665_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_665_select = {
                             in_data[663],
                             in_data[182],
                             in_data[27],
                             in_data[168],
                             in_data[399],
                             in_data[31]};
    
    wire lut_665_out = lut_665_table[lut_665_select];
    
    generate
    if ( USE_REG ) begin : ff_665
        reg   lut_665_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_665_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_665_ff <= lut_665_out;
            end
        end
        
        assign out_data[665] = lut_665_ff;
    end
    else begin : no_ff_665
        assign out_data[665] = lut_665_out;
    end
    endgenerate
    
    
    
    // LUT : 666
    wire [63:0] lut_666_table = 64'b0000000000000000001000100010001000000000000000001011101110111011;
    wire [5:0] lut_666_select = {
                             in_data[314],
                             in_data[579],
                             in_data[254],
                             in_data[503],
                             in_data[287],
                             in_data[407]};
    
    wire lut_666_out = lut_666_table[lut_666_select];
    
    generate
    if ( USE_REG ) begin : ff_666
        reg   lut_666_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_666_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_666_ff <= lut_666_out;
            end
        end
        
        assign out_data[666] = lut_666_ff;
    end
    else begin : no_ff_666
        assign out_data[666] = lut_666_out;
    end
    endgenerate
    
    
    
    // LUT : 667
    wire [63:0] lut_667_table = 64'b0000000000000000000011000000000000001111001111110100110011111111;
    wire [5:0] lut_667_select = {
                             in_data[239],
                             in_data[426],
                             in_data[609],
                             in_data[570],
                             in_data[351],
                             in_data[588]};
    
    wire lut_667_out = lut_667_table[lut_667_select];
    
    generate
    if ( USE_REG ) begin : ff_667
        reg   lut_667_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_667_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_667_ff <= lut_667_out;
            end
        end
        
        assign out_data[667] = lut_667_ff;
    end
    else begin : no_ff_667
        assign out_data[667] = lut_667_out;
    end
    endgenerate
    
    
    
    // LUT : 668
    wire [63:0] lut_668_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_668_select = {
                             in_data[289],
                             in_data[139],
                             in_data[771],
                             in_data[0],
                             in_data[685],
                             in_data[750]};
    
    wire lut_668_out = lut_668_table[lut_668_select];
    
    generate
    if ( USE_REG ) begin : ff_668
        reg   lut_668_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_668_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_668_ff <= lut_668_out;
            end
        end
        
        assign out_data[668] = lut_668_ff;
    end
    else begin : no_ff_668
        assign out_data[668] = lut_668_out;
    end
    endgenerate
    
    
    
    // LUT : 669
    wire [63:0] lut_669_table = 64'b1111111110101010111111111000101011111111000010101111111100000000;
    wire [5:0] lut_669_select = {
                             in_data[521],
                             in_data[623],
                             in_data[159],
                             in_data[740],
                             in_data[76],
                             in_data[405]};
    
    wire lut_669_out = lut_669_table[lut_669_select];
    
    generate
    if ( USE_REG ) begin : ff_669
        reg   lut_669_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_669_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_669_ff <= lut_669_out;
            end
        end
        
        assign out_data[669] = lut_669_ff;
    end
    else begin : no_ff_669
        assign out_data[669] = lut_669_out;
    end
    endgenerate
    
    
    
    // LUT : 670
    wire [63:0] lut_670_table = 64'b0000000000110011000000000011001100000000001100110000000000110011;
    wire [5:0] lut_670_select = {
                             in_data[774],
                             in_data[699],
                             in_data[569],
                             in_data[334],
                             in_data[360],
                             in_data[74]};
    
    wire lut_670_out = lut_670_table[lut_670_select];
    
    generate
    if ( USE_REG ) begin : ff_670
        reg   lut_670_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_670_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_670_ff <= lut_670_out;
            end
        end
        
        assign out_data[670] = lut_670_ff;
    end
    else begin : no_ff_670
        assign out_data[670] = lut_670_out;
    end
    endgenerate
    
    
    
    // LUT : 671
    wire [63:0] lut_671_table = 64'b0001111100001111000001010000010100011111000011110000110100000101;
    wire [5:0] lut_671_select = {
                             in_data[250],
                             in_data[359],
                             in_data[80],
                             in_data[630],
                             in_data[170],
                             in_data[259]};
    
    wire lut_671_out = lut_671_table[lut_671_select];
    
    generate
    if ( USE_REG ) begin : ff_671
        reg   lut_671_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_671_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_671_ff <= lut_671_out;
            end
        end
        
        assign out_data[671] = lut_671_ff;
    end
    else begin : no_ff_671
        assign out_data[671] = lut_671_out;
    end
    endgenerate
    
    
    
    // LUT : 672
    wire [63:0] lut_672_table = 64'b0000000000000001000000000000000100000001000000010000000100000001;
    wire [5:0] lut_672_select = {
                             in_data[269],
                             in_data[82],
                             in_data[756],
                             in_data[566],
                             in_data[332],
                             in_data[161]};
    
    wire lut_672_out = lut_672_table[lut_672_select];
    
    generate
    if ( USE_REG ) begin : ff_672
        reg   lut_672_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_672_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_672_ff <= lut_672_out;
            end
        end
        
        assign out_data[672] = lut_672_ff;
    end
    else begin : no_ff_672
        assign out_data[672] = lut_672_out;
    end
    endgenerate
    
    
    
    // LUT : 673
    wire [63:0] lut_673_table = 64'b1111111111111111111111110000000011111111111111111111111100000000;
    wire [5:0] lut_673_select = {
                             in_data[615],
                             in_data[209],
                             in_data[451],
                             in_data[747],
                             in_data[729],
                             in_data[419]};
    
    wire lut_673_out = lut_673_table[lut_673_select];
    
    generate
    if ( USE_REG ) begin : ff_673
        reg   lut_673_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_673_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_673_ff <= lut_673_out;
            end
        end
        
        assign out_data[673] = lut_673_ff;
    end
    else begin : no_ff_673
        assign out_data[673] = lut_673_out;
    end
    endgenerate
    
    
    
    // LUT : 674
    wire [63:0] lut_674_table = 64'b1111111111111111111111111111111110001011000000100000111100000010;
    wire [5:0] lut_674_select = {
                             in_data[539],
                             in_data[767],
                             in_data[660],
                             in_data[574],
                             in_data[175],
                             in_data[236]};
    
    wire lut_674_out = lut_674_table[lut_674_select];
    
    generate
    if ( USE_REG ) begin : ff_674
        reg   lut_674_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_674_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_674_ff <= lut_674_out;
            end
        end
        
        assign out_data[674] = lut_674_ff;
    end
    else begin : no_ff_674
        assign out_data[674] = lut_674_out;
    end
    endgenerate
    
    
    
    // LUT : 675
    wire [63:0] lut_675_table = 64'b1111111111111111000000000000000011111111111111110000111100001111;
    wire [5:0] lut_675_select = {
                             in_data[458],
                             in_data[689],
                             in_data[64],
                             in_data[434],
                             in_data[646],
                             in_data[578]};
    
    wire lut_675_out = lut_675_table[lut_675_select];
    
    generate
    if ( USE_REG ) begin : ff_675
        reg   lut_675_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_675_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_675_ff <= lut_675_out;
            end
        end
        
        assign out_data[675] = lut_675_ff;
    end
    else begin : no_ff_675
        assign out_data[675] = lut_675_out;
    end
    endgenerate
    
    
    
    // LUT : 676
    wire [63:0] lut_676_table = 64'b1101110101010101110111010101010111011101010101011101110101010101;
    wire [5:0] lut_676_select = {
                             in_data[704],
                             in_data[697],
                             in_data[542],
                             in_data[590],
                             in_data[123],
                             in_data[375]};
    
    wire lut_676_out = lut_676_table[lut_676_select];
    
    generate
    if ( USE_REG ) begin : ff_676
        reg   lut_676_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_676_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_676_ff <= lut_676_out;
            end
        end
        
        assign out_data[676] = lut_676_ff;
    end
    else begin : no_ff_676
        assign out_data[676] = lut_676_out;
    end
    endgenerate
    
    
    
    // LUT : 677
    wire [63:0] lut_677_table = 64'b0000000011101110101000001111111010101010111111101010101011111110;
    wire [5:0] lut_677_select = {
                             in_data[44],
                             in_data[144],
                             in_data[156],
                             in_data[640],
                             in_data[438],
                             in_data[716]};
    
    wire lut_677_out = lut_677_table[lut_677_select];
    
    generate
    if ( USE_REG ) begin : ff_677
        reg   lut_677_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_677_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_677_ff <= lut_677_out;
            end
        end
        
        assign out_data[677] = lut_677_ff;
    end
    else begin : no_ff_677
        assign out_data[677] = lut_677_out;
    end
    endgenerate
    
    
    
    // LUT : 678
    wire [63:0] lut_678_table = 64'b0000010000000000000001000000010000000101000001010000010100000101;
    wire [5:0] lut_678_select = {
                             in_data[772],
                             in_data[51],
                             in_data[143],
                             in_data[317],
                             in_data[506],
                             in_data[340]};
    
    wire lut_678_out = lut_678_table[lut_678_select];
    
    generate
    if ( USE_REG ) begin : ff_678
        reg   lut_678_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_678_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_678_ff <= lut_678_out;
            end
        end
        
        assign out_data[678] = lut_678_ff;
    end
    else begin : no_ff_678
        assign out_data[678] = lut_678_out;
    end
    endgenerate
    
    
    
    // LUT : 679
    wire [63:0] lut_679_table = 64'b1111111111111111000001010000000011111111111111110011101100000000;
    wire [5:0] lut_679_select = {
                             in_data[169],
                             in_data[576],
                             in_data[52],
                             in_data[477],
                             in_data[33],
                             in_data[761]};
    
    wire lut_679_out = lut_679_table[lut_679_select];
    
    generate
    if ( USE_REG ) begin : ff_679
        reg   lut_679_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_679_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_679_ff <= lut_679_out;
            end
        end
        
        assign out_data[679] = lut_679_ff;
    end
    else begin : no_ff_679
        assign out_data[679] = lut_679_out;
    end
    endgenerate
    
    
    
    // LUT : 680
    wire [63:0] lut_680_table = 64'b1010111111111111000000000000101010100111111111110000000000000000;
    wire [5:0] lut_680_select = {
                             in_data[418],
                             in_data[550],
                             in_data[202],
                             in_data[564],
                             in_data[769],
                             in_data[207]};
    
    wire lut_680_out = lut_680_table[lut_680_select];
    
    generate
    if ( USE_REG ) begin : ff_680
        reg   lut_680_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_680_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_680_ff <= lut_680_out;
            end
        end
        
        assign out_data[680] = lut_680_ff;
    end
    else begin : no_ff_680
        assign out_data[680] = lut_680_out;
    end
    endgenerate
    
    
    
    // LUT : 681
    wire [63:0] lut_681_table = 64'b0000000000010001000000000000000000000000101111110000000010101111;
    wire [5:0] lut_681_select = {
                             in_data[627],
                             in_data[273],
                             in_data[147],
                             in_data[179],
                             in_data[111],
                             in_data[691]};
    
    wire lut_681_out = lut_681_table[lut_681_select];
    
    generate
    if ( USE_REG ) begin : ff_681
        reg   lut_681_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_681_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_681_ff <= lut_681_out;
            end
        end
        
        assign out_data[681] = lut_681_ff;
    end
    else begin : no_ff_681
        assign out_data[681] = lut_681_out;
    end
    endgenerate
    
    
    
    // LUT : 682
    wire [63:0] lut_682_table = 64'b0000000001010001000100010101000100010011010101010001001101010101;
    wire [5:0] lut_682_select = {
                             in_data[748],
                             in_data[727],
                             in_data[469],
                             in_data[215],
                             in_data[343],
                             in_data[324]};
    
    wire lut_682_out = lut_682_table[lut_682_select];
    
    generate
    if ( USE_REG ) begin : ff_682
        reg   lut_682_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_682_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_682_ff <= lut_682_out;
            end
        end
        
        assign out_data[682] = lut_682_ff;
    end
    else begin : no_ff_682
        assign out_data[682] = lut_682_out;
    end
    endgenerate
    
    
    
    // LUT : 683
    wire [63:0] lut_683_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_683_select = {
                             in_data[37],
                             in_data[53],
                             in_data[246],
                             in_data[768],
                             in_data[140],
                             in_data[679]};
    
    wire lut_683_out = lut_683_table[lut_683_select];
    
    generate
    if ( USE_REG ) begin : ff_683
        reg   lut_683_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_683_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_683_ff <= lut_683_out;
            end
        end
        
        assign out_data[683] = lut_683_ff;
    end
    else begin : no_ff_683
        assign out_data[683] = lut_683_out;
    end
    endgenerate
    
    
    
    // LUT : 684
    wire [63:0] lut_684_table = 64'b0101010101010101010101010100000001110101010101010101010101000000;
    wire [5:0] lut_684_select = {
                             in_data[196],
                             in_data[459],
                             in_data[629],
                             in_data[303],
                             in_data[228],
                             in_data[356]};
    
    wire lut_684_out = lut_684_table[lut_684_select];
    
    generate
    if ( USE_REG ) begin : ff_684
        reg   lut_684_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_684_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_684_ff <= lut_684_out;
            end
        end
        
        assign out_data[684] = lut_684_ff;
    end
    else begin : no_ff_684
        assign out_data[684] = lut_684_out;
    end
    endgenerate
    
    
    
    // LUT : 685
    wire [63:0] lut_685_table = 64'b1111111111111011101100111011001011110111111110111011001010100010;
    wire [5:0] lut_685_select = {
                             in_data[187],
                             in_data[555],
                             in_data[462],
                             in_data[567],
                             in_data[105],
                             in_data[398]};
    
    wire lut_685_out = lut_685_table[lut_685_select];
    
    generate
    if ( USE_REG ) begin : ff_685
        reg   lut_685_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_685_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_685_ff <= lut_685_out;
            end
        end
        
        assign out_data[685] = lut_685_ff;
    end
    else begin : no_ff_685
        assign out_data[685] = lut_685_out;
    end
    endgenerate
    
    
    
    // LUT : 686
    wire [63:0] lut_686_table = 64'b0000000000000000000000000000000010101010001010101010101110101111;
    wire [5:0] lut_686_select = {
                             in_data[491],
                             in_data[723],
                             in_data[502],
                             in_data[667],
                             in_data[79],
                             in_data[676]};
    
    wire lut_686_out = lut_686_table[lut_686_select];
    
    generate
    if ( USE_REG ) begin : ff_686
        reg   lut_686_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_686_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_686_ff <= lut_686_out;
            end
        end
        
        assign out_data[686] = lut_686_ff;
    end
    else begin : no_ff_686
        assign out_data[686] = lut_686_out;
    end
    endgenerate
    
    
    
    // LUT : 687
    wire [63:0] lut_687_table = 64'b1110111000000000111111110000000011111111000000011111111100000000;
    wire [5:0] lut_687_select = {
                             in_data[732],
                             in_data[21],
                             in_data[406],
                             in_data[253],
                             in_data[738],
                             in_data[258]};
    
    wire lut_687_out = lut_687_table[lut_687_select];
    
    generate
    if ( USE_REG ) begin : ff_687
        reg   lut_687_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_687_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_687_ff <= lut_687_out;
            end
        end
        
        assign out_data[687] = lut_687_ff;
    end
    else begin : no_ff_687
        assign out_data[687] = lut_687_out;
    end
    endgenerate
    
    
    
    // LUT : 688
    wire [63:0] lut_688_table = 64'b1011101110111011100110101001101010111011101110111011101010011010;
    wire [5:0] lut_688_select = {
                             in_data[9],
                             in_data[528],
                             in_data[562],
                             in_data[220],
                             in_data[572],
                             in_data[514]};
    
    wire lut_688_out = lut_688_table[lut_688_select];
    
    generate
    if ( USE_REG ) begin : ff_688
        reg   lut_688_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_688_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_688_ff <= lut_688_out;
            end
        end
        
        assign out_data[688] = lut_688_ff;
    end
    else begin : no_ff_688
        assign out_data[688] = lut_688_out;
    end
    endgenerate
    
    
    
    // LUT : 689
    wire [63:0] lut_689_table = 64'b1010101010101010101110111010101010101010101010101011101110101010;
    wire [5:0] lut_689_select = {
                             in_data[632],
                             in_data[77],
                             in_data[613],
                             in_data[450],
                             in_data[70],
                             in_data[229]};
    
    wire lut_689_out = lut_689_table[lut_689_select];
    
    generate
    if ( USE_REG ) begin : ff_689
        reg   lut_689_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_689_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_689_ff <= lut_689_out;
            end
        end
        
        assign out_data[689] = lut_689_ff;
    end
    else begin : no_ff_689
        assign out_data[689] = lut_689_out;
    end
    endgenerate
    
    
    
    // LUT : 690
    wire [63:0] lut_690_table = 64'b0000000000000000111111111101110100000000000000001111111101011101;
    wire [5:0] lut_690_select = {
                             in_data[775],
                             in_data[271],
                             in_data[176],
                             in_data[63],
                             in_data[776],
                             in_data[305]};
    
    wire lut_690_out = lut_690_table[lut_690_select];
    
    generate
    if ( USE_REG ) begin : ff_690
        reg   lut_690_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_690_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_690_ff <= lut_690_out;
            end
        end
        
        assign out_data[690] = lut_690_ff;
    end
    else begin : no_ff_690
        assign out_data[690] = lut_690_out;
    end
    endgenerate
    
    
    
    // LUT : 691
    wire [63:0] lut_691_table = 64'b0011001100110011001100110001001100110011000100110001001100010011;
    wire [5:0] lut_691_select = {
                             in_data[40],
                             in_data[643],
                             in_data[107],
                             in_data[181],
                             in_data[551],
                             in_data[242]};
    
    wire lut_691_out = lut_691_table[lut_691_select];
    
    generate
    if ( USE_REG ) begin : ff_691
        reg   lut_691_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_691_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_691_ff <= lut_691_out;
            end
        end
        
        assign out_data[691] = lut_691_ff;
    end
    else begin : no_ff_691
        assign out_data[691] = lut_691_out;
    end
    endgenerate
    
    
    
    // LUT : 692
    wire [63:0] lut_692_table = 64'b0111010000000000000000000000000011111111111111110000000011111111;
    wire [5:0] lut_692_select = {
                             in_data[461],
                             in_data[626],
                             in_data[155],
                             in_data[3],
                             in_data[2],
                             in_data[59]};
    
    wire lut_692_out = lut_692_table[lut_692_select];
    
    generate
    if ( USE_REG ) begin : ff_692
        reg   lut_692_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_692_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_692_ff <= lut_692_out;
            end
        end
        
        assign out_data[692] = lut_692_ff;
    end
    else begin : no_ff_692
        assign out_data[692] = lut_692_out;
    end
    endgenerate
    
    
    
    // LUT : 693
    wire [63:0] lut_693_table = 64'b1111011111111111111100001111110011111111111111110000000011111100;
    wire [5:0] lut_693_select = {
                             in_data[400],
                             in_data[150],
                             in_data[153],
                             in_data[104],
                             in_data[624],
                             in_data[672]};
    
    wire lut_693_out = lut_693_table[lut_693_select];
    
    generate
    if ( USE_REG ) begin : ff_693
        reg   lut_693_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_693_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_693_ff <= lut_693_out;
            end
        end
        
        assign out_data[693] = lut_693_ff;
    end
    else begin : no_ff_693
        assign out_data[693] = lut_693_out;
    end
    endgenerate
    
    
    
    // LUT : 694
    wire [63:0] lut_694_table = 64'b0000000000000000111111110011001100000000000000000000001100000011;
    wire [5:0] lut_694_select = {
                             in_data[439],
                             in_data[719],
                             in_data[648],
                             in_data[659],
                             in_data[186],
                             in_data[535]};
    
    wire lut_694_out = lut_694_table[lut_694_select];
    
    generate
    if ( USE_REG ) begin : ff_694
        reg   lut_694_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_694_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_694_ff <= lut_694_out;
            end
        end
        
        assign out_data[694] = lut_694_ff;
    end
    else begin : no_ff_694
        assign out_data[694] = lut_694_out;
    end
    endgenerate
    
    
    
    // LUT : 695
    wire [63:0] lut_695_table = 64'b0011011100110111001101110011011101110101011101010111010101110111;
    wire [5:0] lut_695_select = {
                             in_data[428],
                             in_data[753],
                             in_data[57],
                             in_data[238],
                             in_data[212],
                             in_data[601]};
    
    wire lut_695_out = lut_695_table[lut_695_select];
    
    generate
    if ( USE_REG ) begin : ff_695
        reg   lut_695_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_695_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_695_ff <= lut_695_out;
            end
        end
        
        assign out_data[695] = lut_695_ff;
    end
    else begin : no_ff_695
        assign out_data[695] = lut_695_out;
    end
    endgenerate
    
    
    
    // LUT : 696
    wire [63:0] lut_696_table = 64'b0001010100010101000000010000000100010101000101010000000100000001;
    wire [5:0] lut_696_select = {
                             in_data[114],
                             in_data[389],
                             in_data[224],
                             in_data[654],
                             in_data[135],
                             in_data[276]};
    
    wire lut_696_out = lut_696_table[lut_696_select];
    
    generate
    if ( USE_REG ) begin : ff_696
        reg   lut_696_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_696_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_696_ff <= lut_696_out;
            end
        end
        
        assign out_data[696] = lut_696_ff;
    end
    else begin : no_ff_696
        assign out_data[696] = lut_696_out;
    end
    endgenerate
    
    
    
    // LUT : 697
    wire [63:0] lut_697_table = 64'b1111111111111111111111111111111111111111111111111101000011010000;
    wire [5:0] lut_697_select = {
                             in_data[412],
                             in_data[425],
                             in_data[5],
                             in_data[71],
                             in_data[733],
                             in_data[120]};
    
    wire lut_697_out = lut_697_table[lut_697_select];
    
    generate
    if ( USE_REG ) begin : ff_697
        reg   lut_697_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_697_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_697_ff <= lut_697_out;
            end
        end
        
        assign out_data[697] = lut_697_ff;
    end
    else begin : no_ff_697
        assign out_data[697] = lut_697_out;
    end
    endgenerate
    
    
    
    // LUT : 698
    wire [63:0] lut_698_table = 64'b0000000000000000000000000100110000000000010011001100110011111111;
    wire [5:0] lut_698_select = {
                             in_data[483],
                             in_data[721],
                             in_data[65],
                             in_data[113],
                             in_data[658],
                             in_data[162]};
    
    wire lut_698_out = lut_698_table[lut_698_select];
    
    generate
    if ( USE_REG ) begin : ff_698
        reg   lut_698_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_698_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_698_ff <= lut_698_out;
            end
        end
        
        assign out_data[698] = lut_698_ff;
    end
    else begin : no_ff_698
        assign out_data[698] = lut_698_out;
    end
    endgenerate
    
    
    
    // LUT : 699
    wire [63:0] lut_699_table = 64'b1110111110001100110111111100110011111111110011001111111111001100;
    wire [5:0] lut_699_select = {
                             in_data[696],
                             in_data[645],
                             in_data[148],
                             in_data[142],
                             in_data[499],
                             in_data[364]};
    
    wire lut_699_out = lut_699_table[lut_699_select];
    
    generate
    if ( USE_REG ) begin : ff_699
        reg   lut_699_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_699_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_699_ff <= lut_699_out;
            end
        end
        
        assign out_data[699] = lut_699_ff;
    end
    else begin : no_ff_699
        assign out_data[699] = lut_699_out;
    end
    endgenerate
    
    
    
    // LUT : 700
    wire [63:0] lut_700_table = 64'b1111101111111111111110111111111100100000101100110010000010110011;
    wire [5:0] lut_700_select = {
                             in_data[444],
                             in_data[702],
                             in_data[424],
                             in_data[669],
                             in_data[372],
                             in_data[174]};
    
    wire lut_700_out = lut_700_table[lut_700_select];
    
    generate
    if ( USE_REG ) begin : ff_700
        reg   lut_700_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_700_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_700_ff <= lut_700_out;
            end
        end
        
        assign out_data[700] = lut_700_ff;
    end
    else begin : no_ff_700
        assign out_data[700] = lut_700_out;
    end
    endgenerate
    
    
    
    // LUT : 701
    wire [63:0] lut_701_table = 64'b1101000011010000111101001111010001010000010101011101010101000100;
    wire [5:0] lut_701_select = {
                             in_data[602],
                             in_data[415],
                             in_data[39],
                             in_data[628],
                             in_data[201],
                             in_data[68]};
    
    wire lut_701_out = lut_701_table[lut_701_select];
    
    generate
    if ( USE_REG ) begin : ff_701
        reg   lut_701_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_701_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_701_ff <= lut_701_out;
            end
        end
        
        assign out_data[701] = lut_701_ff;
    end
    else begin : no_ff_701
        assign out_data[701] = lut_701_out;
    end
    endgenerate
    
    
    
    // LUT : 702
    wire [63:0] lut_702_table = 64'b0000000011001100000000001101111100000000111111110000000011111111;
    wire [5:0] lut_702_select = {
                             in_data[296],
                             in_data[252],
                             in_data[320],
                             in_data[448],
                             in_data[95],
                             in_data[141]};
    
    wire lut_702_out = lut_702_table[lut_702_select];
    
    generate
    if ( USE_REG ) begin : ff_702
        reg   lut_702_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_702_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_702_ff <= lut_702_out;
            end
        end
        
        assign out_data[702] = lut_702_ff;
    end
    else begin : no_ff_702
        assign out_data[702] = lut_702_out;
    end
    endgenerate
    
    
    
    // LUT : 703
    wire [63:0] lut_703_table = 64'b1111111110101111001000101010001000100010101000100010101010101010;
    wire [5:0] lut_703_select = {
                             in_data[525],
                             in_data[342],
                             in_data[341],
                             in_data[377],
                             in_data[687],
                             in_data[378]};
    
    wire lut_703_out = lut_703_table[lut_703_select];
    
    generate
    if ( USE_REG ) begin : ff_703
        reg   lut_703_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_703_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_703_ff <= lut_703_out;
            end
        end
        
        assign out_data[703] = lut_703_ff;
    end
    else begin : no_ff_703
        assign out_data[703] = lut_703_out;
    end
    endgenerate
    
    
    
    // LUT : 704
    wire [63:0] lut_704_table = 64'b1111111100001011111111110000111111111111000010111011111100001111;
    wire [5:0] lut_704_select = {
                             in_data[199],
                             in_data[442],
                             in_data[369],
                             in_data[291],
                             in_data[98],
                             in_data[128]};
    
    wire lut_704_out = lut_704_table[lut_704_select];
    
    generate
    if ( USE_REG ) begin : ff_704
        reg   lut_704_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_704_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_704_ff <= lut_704_out;
            end
        end
        
        assign out_data[704] = lut_704_ff;
    end
    else begin : no_ff_704
        assign out_data[704] = lut_704_out;
    end
    endgenerate
    
    
    
    // LUT : 705
    wire [63:0] lut_705_table = 64'b1111001111111111111100111111111111110000111100111111000011110011;
    wire [5:0] lut_705_select = {
                             in_data[72],
                             in_data[11],
                             in_data[339],
                             in_data[472],
                             in_data[180],
                             in_data[14]};
    
    wire lut_705_out = lut_705_table[lut_705_select];
    
    generate
    if ( USE_REG ) begin : ff_705
        reg   lut_705_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_705_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_705_ff <= lut_705_out;
            end
        end
        
        assign out_data[705] = lut_705_ff;
    end
    else begin : no_ff_705
        assign out_data[705] = lut_705_out;
    end
    endgenerate
    
    
    
    // LUT : 706
    wire [63:0] lut_706_table = 64'b1111111110100000111111110000100011111111001100001111111100110011;
    wire [5:0] lut_706_select = {
                             in_data[457],
                             in_data[330],
                             in_data[594],
                             in_data[383],
                             in_data[430],
                             in_data[23]};
    
    wire lut_706_out = lut_706_table[lut_706_select];
    
    generate
    if ( USE_REG ) begin : ff_706
        reg   lut_706_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_706_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_706_ff <= lut_706_out;
            end
        end
        
        assign out_data[706] = lut_706_ff;
    end
    else begin : no_ff_706
        assign out_data[706] = lut_706_out;
    end
    endgenerate
    
    
    
    // LUT : 707
    wire [63:0] lut_707_table = 64'b1101110111111111111111111111111111010000110100011010000010101010;
    wire [5:0] lut_707_select = {
                             in_data[152],
                             in_data[189],
                             in_data[423],
                             in_data[92],
                             in_data[527],
                             in_data[268]};
    
    wire lut_707_out = lut_707_table[lut_707_select];
    
    generate
    if ( USE_REG ) begin : ff_707
        reg   lut_707_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_707_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_707_ff <= lut_707_out;
            end
        end
        
        assign out_data[707] = lut_707_ff;
    end
    else begin : no_ff_707
        assign out_data[707] = lut_707_out;
    end
    endgenerate
    
    
    
    // LUT : 708
    wire [63:0] lut_708_table = 64'b0000000011111111001100000010001100000000111111110011000000000011;
    wire [5:0] lut_708_select = {
                             in_data[15],
                             in_data[636],
                             in_data[599],
                             in_data[519],
                             in_data[286],
                             in_data[367]};
    
    wire lut_708_out = lut_708_table[lut_708_select];
    
    generate
    if ( USE_REG ) begin : ff_708
        reg   lut_708_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_708_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_708_ff <= lut_708_out;
            end
        end
        
        assign out_data[708] = lut_708_ff;
    end
    else begin : no_ff_708
        assign out_data[708] = lut_708_out;
    end
    endgenerate
    
    
    
    // LUT : 709
    wire [63:0] lut_709_table = 64'b0011000000110000001100110011000000110000001100000011000100110000;
    wire [5:0] lut_709_select = {
                             in_data[43],
                             in_data[119],
                             in_data[49],
                             in_data[157],
                             in_data[664],
                             in_data[54]};
    
    wire lut_709_out = lut_709_table[lut_709_select];
    
    generate
    if ( USE_REG ) begin : ff_709
        reg   lut_709_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_709_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_709_ff <= lut_709_out;
            end
        end
        
        assign out_data[709] = lut_709_ff;
    end
    else begin : no_ff_709
        assign out_data[709] = lut_709_out;
    end
    endgenerate
    
    
    
    // LUT : 710
    wire [63:0] lut_710_table = 64'b0000000000000000000000000000000000010001000100010000001100010011;
    wire [5:0] lut_710_select = {
                             in_data[132],
                             in_data[610],
                             in_data[282],
                             in_data[311],
                             in_data[711],
                             in_data[635]};
    
    wire lut_710_out = lut_710_table[lut_710_select];
    
    generate
    if ( USE_REG ) begin : ff_710
        reg   lut_710_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_710_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_710_ff <= lut_710_out;
            end
        end
        
        assign out_data[710] = lut_710_ff;
    end
    else begin : no_ff_710
        assign out_data[710] = lut_710_out;
    end
    endgenerate
    
    
    
    // LUT : 711
    wire [63:0] lut_711_table = 64'b1100111111001111000011110000111111001111110011110000111100001101;
    wire [5:0] lut_711_select = {
                             in_data[30],
                             in_data[158],
                             in_data[600],
                             in_data[522],
                             in_data[354],
                             in_data[112]};
    
    wire lut_711_out = lut_711_table[lut_711_select];
    
    generate
    if ( USE_REG ) begin : ff_711
        reg   lut_711_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_711_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_711_ff <= lut_711_out;
            end
        end
        
        assign out_data[711] = lut_711_ff;
    end
    else begin : no_ff_711
        assign out_data[711] = lut_711_out;
    end
    endgenerate
    
    
    
    // LUT : 712
    wire [63:0] lut_712_table = 64'b0111011100110111000000000011000101111111001101110000000000110011;
    wire [5:0] lut_712_select = {
                             in_data[47],
                             in_data[651],
                             in_data[403],
                             in_data[587],
                             in_data[134],
                             in_data[164]};
    
    wire lut_712_out = lut_712_table[lut_712_select];
    
    generate
    if ( USE_REG ) begin : ff_712
        reg   lut_712_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_712_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_712_ff <= lut_712_out;
            end
        end
        
        assign out_data[712] = lut_712_ff;
    end
    else begin : no_ff_712
        assign out_data[712] = lut_712_out;
    end
    endgenerate
    
    
    
    // LUT : 713
    wire [63:0] lut_713_table = 64'b0000000011011100000000000101000001000000110111010001000001110001;
    wire [5:0] lut_713_select = {
                             in_data[481],
                             in_data[580],
                             in_data[453],
                             in_data[577],
                             in_data[414],
                             in_data[486]};
    
    wire lut_713_out = lut_713_table[lut_713_select];
    
    generate
    if ( USE_REG ) begin : ff_713
        reg   lut_713_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_713_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_713_ff <= lut_713_out;
            end
        end
        
        assign out_data[713] = lut_713_ff;
    end
    else begin : no_ff_713
        assign out_data[713] = lut_713_out;
    end
    endgenerate
    
    
    
    // LUT : 714
    wire [63:0] lut_714_table = 64'b0101010101110101010101010111010101110101011101010111000101110101;
    wire [5:0] lut_714_select = {
                             in_data[353],
                             in_data[730],
                             in_data[598],
                             in_data[409],
                             in_data[355],
                             in_data[241]};
    
    wire lut_714_out = lut_714_table[lut_714_select];
    
    generate
    if ( USE_REG ) begin : ff_714
        reg   lut_714_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_714_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_714_ff <= lut_714_out;
            end
        end
        
        assign out_data[714] = lut_714_ff;
    end
    else begin : no_ff_714
        assign out_data[714] = lut_714_out;
    end
    endgenerate
    
    
    
    // LUT : 715
    wire [63:0] lut_715_table = 64'b0010001000100010111100100011001011101111101011111111111111111111;
    wire [5:0] lut_715_select = {
                             in_data[185],
                             in_data[489],
                             in_data[85],
                             in_data[243],
                             in_data[410],
                             in_data[387]};
    
    wire lut_715_out = lut_715_table[lut_715_select];
    
    generate
    if ( USE_REG ) begin : ff_715
        reg   lut_715_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_715_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_715_ff <= lut_715_out;
            end
        end
        
        assign out_data[715] = lut_715_ff;
    end
    else begin : no_ff_715
        assign out_data[715] = lut_715_out;
    end
    endgenerate
    
    
    
    // LUT : 716
    wire [63:0] lut_716_table = 64'b1111111111111111111111011111111111110100111111110001000011111111;
    wire [5:0] lut_716_select = {
                             in_data[284],
                             in_data[255],
                             in_data[402],
                             in_data[737],
                             in_data[365],
                             in_data[106]};
    
    wire lut_716_out = lut_716_table[lut_716_select];
    
    generate
    if ( USE_REG ) begin : ff_716
        reg   lut_716_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_716_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_716_ff <= lut_716_out;
            end
        end
        
        assign out_data[716] = lut_716_ff;
    end
    else begin : no_ff_716
        assign out_data[716] = lut_716_out;
    end
    endgenerate
    
    
    
    // LUT : 717
    wire [63:0] lut_717_table = 64'b0000000000100010000000000011001100000000000000000000000000110011;
    wire [5:0] lut_717_select = {
                             in_data[653],
                             in_data[739],
                             in_data[515],
                             in_data[223],
                             in_data[556],
                             in_data[455]};
    
    wire lut_717_out = lut_717_table[lut_717_select];
    
    generate
    if ( USE_REG ) begin : ff_717
        reg   lut_717_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_717_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_717_ff <= lut_717_out;
            end
        end
        
        assign out_data[717] = lut_717_ff;
    end
    else begin : no_ff_717
        assign out_data[717] = lut_717_out;
    end
    endgenerate
    
    
    
    // LUT : 718
    wire [63:0] lut_718_table = 64'b0000111111111111111100011111000001011111010101011111010111110000;
    wire [5:0] lut_718_select = {
                             in_data[101],
                             in_data[662],
                             in_data[208],
                             in_data[244],
                             in_data[504],
                             in_data[668]};
    
    wire lut_718_out = lut_718_table[lut_718_select];
    
    generate
    if ( USE_REG ) begin : ff_718
        reg   lut_718_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_718_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_718_ff <= lut_718_out;
            end
        end
        
        assign out_data[718] = lut_718_ff;
    end
    else begin : no_ff_718
        assign out_data[718] = lut_718_out;
    end
    endgenerate
    
    
    
    // LUT : 719
    wire [63:0] lut_719_table = 64'b1111111111111111111111111111101011111111111111111111101011111010;
    wire [5:0] lut_719_select = {
                             in_data[682],
                             in_data[688],
                             in_data[540],
                             in_data[583],
                             in_data[16],
                             in_data[302]};
    
    wire lut_719_out = lut_719_table[lut_719_select];
    
    generate
    if ( USE_REG ) begin : ff_719
        reg   lut_719_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_719_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_719_ff <= lut_719_out;
            end
        end
        
        assign out_data[719] = lut_719_ff;
    end
    else begin : no_ff_719
        assign out_data[719] = lut_719_out;
    end
    endgenerate
    
    
    
    // LUT : 720
    wire [63:0] lut_720_table = 64'b0000000011110011000000000111001100000000111100110000000011110011;
    wire [5:0] lut_720_select = {
                             in_data[29],
                             in_data[530],
                             in_data[652],
                             in_data[136],
                             in_data[206],
                             in_data[22]};
    
    wire lut_720_out = lut_720_table[lut_720_select];
    
    generate
    if ( USE_REG ) begin : ff_720
        reg   lut_720_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_720_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_720_ff <= lut_720_out;
            end
        end
        
        assign out_data[720] = lut_720_ff;
    end
    else begin : no_ff_720
        assign out_data[720] = lut_720_out;
    end
    endgenerate
    
    
    
    // LUT : 721
    wire [63:0] lut_721_table = 64'b1010101011111111101010101111111110101010111111111010101011111111;
    wire [5:0] lut_721_select = {
                             in_data[12],
                             in_data[171],
                             in_data[440],
                             in_data[281],
                             in_data[357],
                             in_data[720]};
    
    wire lut_721_out = lut_721_table[lut_721_select];
    
    generate
    if ( USE_REG ) begin : ff_721
        reg   lut_721_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_721_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_721_ff <= lut_721_out;
            end
        end
        
        assign out_data[721] = lut_721_ff;
    end
    else begin : no_ff_721
        assign out_data[721] = lut_721_out;
    end
    endgenerate
    
    
    
    // LUT : 722
    wire [63:0] lut_722_table = 64'b0000000000001010000000000101111100000000000010100000000000011111;
    wire [5:0] lut_722_select = {
                             in_data[118],
                             in_data[126],
                             in_data[325],
                             in_data[173],
                             in_data[366],
                             in_data[468]};
    
    wire lut_722_out = lut_722_table[lut_722_select];
    
    generate
    if ( USE_REG ) begin : ff_722
        reg   lut_722_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_722_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_722_ff <= lut_722_out;
            end
        end
        
        assign out_data[722] = lut_722_ff;
    end
    else begin : no_ff_722
        assign out_data[722] = lut_722_out;
    end
    endgenerate
    
    
    
    // LUT : 723
    wire [63:0] lut_723_table = 64'b1110000011100000111000001111000011111110111111001111111011111100;
    wire [5:0] lut_723_select = {
                             in_data[488],
                             in_data[10],
                             in_data[673],
                             in_data[347],
                             in_data[231],
                             in_data[257]};
    
    wire lut_723_out = lut_723_table[lut_723_select];
    
    generate
    if ( USE_REG ) begin : ff_723
        reg   lut_723_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_723_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_723_ff <= lut_723_out;
            end
        end
        
        assign out_data[723] = lut_723_ff;
    end
    else begin : no_ff_723
        assign out_data[723] = lut_723_out;
    end
    endgenerate
    
    
    
    // LUT : 724
    wire [63:0] lut_724_table = 64'b0101000001010000111110101111000011110000111100001111111111111010;
    wire [5:0] lut_724_select = {
                             in_data[557],
                             in_data[445],
                             in_data[219],
                             in_data[686],
                             in_data[394],
                             in_data[348]};
    
    wire lut_724_out = lut_724_table[lut_724_select];
    
    generate
    if ( USE_REG ) begin : ff_724
        reg   lut_724_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_724_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_724_ff <= lut_724_out;
            end
        end
        
        assign out_data[724] = lut_724_ff;
    end
    else begin : no_ff_724
        assign out_data[724] = lut_724_out;
    end
    endgenerate
    
    
    
    // LUT : 725
    wire [63:0] lut_725_table = 64'b0000000000000100100001010000010111000000110001001000000011000100;
    wire [5:0] lut_725_select = {
                             in_data[319],
                             in_data[581],
                             in_data[573],
                             in_data[151],
                             in_data[316],
                             in_data[517]};
    
    wire lut_725_out = lut_725_table[lut_725_select];
    
    generate
    if ( USE_REG ) begin : ff_725
        reg   lut_725_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_725_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_725_ff <= lut_725_out;
            end
        end
        
        assign out_data[725] = lut_725_ff;
    end
    else begin : no_ff_725
        assign out_data[725] = lut_725_out;
    end
    endgenerate
    
    
    
    // LUT : 726
    wire [63:0] lut_726_table = 64'b1010111110101111101011111110111110100000101000001010010010101000;
    wire [5:0] lut_726_select = {
                             in_data[735],
                             in_data[478],
                             in_data[533],
                             in_data[299],
                             in_data[83],
                             in_data[411]};
    
    wire lut_726_out = lut_726_table[lut_726_select];
    
    generate
    if ( USE_REG ) begin : ff_726
        reg   lut_726_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_726_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_726_ff <= lut_726_out;
            end
        end
        
        assign out_data[726] = lut_726_ff;
    end
    else begin : no_ff_726
        assign out_data[726] = lut_726_out;
    end
    endgenerate
    
    
    
    // LUT : 727
    wire [63:0] lut_727_table = 64'b0101110101011111000010000000000001010101010101010000000000000000;
    wire [5:0] lut_727_select = {
                             in_data[338],
                             in_data[379],
                             in_data[266],
                             in_data[500],
                             in_data[310],
                             in_data[358]};
    
    wire lut_727_out = lut_727_table[lut_727_select];
    
    generate
    if ( USE_REG ) begin : ff_727
        reg   lut_727_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_727_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_727_ff <= lut_727_out;
            end
        end
        
        assign out_data[727] = lut_727_ff;
    end
    else begin : no_ff_727
        assign out_data[727] = lut_727_out;
    end
    endgenerate
    
    
    
    // LUT : 728
    wire [63:0] lut_728_table = 64'b1111111111111111111111111111111110110000101100000000000000100000;
    wire [5:0] lut_728_select = {
                             in_data[431],
                             in_data[529],
                             in_data[218],
                             in_data[619],
                             in_data[99],
                             in_data[35]};
    
    wire lut_728_out = lut_728_table[lut_728_select];
    
    generate
    if ( USE_REG ) begin : ff_728
        reg   lut_728_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_728_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_728_ff <= lut_728_out;
            end
        end
        
        assign out_data[728] = lut_728_ff;
    end
    else begin : no_ff_728
        assign out_data[728] = lut_728_out;
    end
    endgenerate
    
    
    
    // LUT : 729
    wire [63:0] lut_729_table = 64'b1111111111111111111111111111111100000000000001000000000000000000;
    wire [5:0] lut_729_select = {
                             in_data[490],
                             in_data[109],
                             in_data[38],
                             in_data[396],
                             in_data[544],
                             in_data[482]};
    
    wire lut_729_out = lut_729_table[lut_729_select];
    
    generate
    if ( USE_REG ) begin : ff_729
        reg   lut_729_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_729_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_729_ff <= lut_729_out;
            end
        end
        
        assign out_data[729] = lut_729_ff;
    end
    else begin : no_ff_729
        assign out_data[729] = lut_729_out;
    end
    endgenerate
    
    
    
    // LUT : 730
    wire [63:0] lut_730_table = 64'b0000000011110011000000001111001100000000111100110000000011110011;
    wire [5:0] lut_730_select = {
                             in_data[392],
                             in_data[87],
                             in_data[596],
                             in_data[712],
                             in_data[270],
                             in_data[703]};
    
    wire lut_730_out = lut_730_table[lut_730_select];
    
    generate
    if ( USE_REG ) begin : ff_730
        reg   lut_730_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_730_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_730_ff <= lut_730_out;
            end
        end
        
        assign out_data[730] = lut_730_ff;
    end
    else begin : no_ff_730
        assign out_data[730] = lut_730_out;
    end
    endgenerate
    
    
    
    // LUT : 731
    wire [63:0] lut_731_table = 64'b0000000011111111000000001111111100000000111011110000000011001111;
    wire [5:0] lut_731_select = {
                             in_data[24],
                             in_data[752],
                             in_data[247],
                             in_data[476],
                             in_data[505],
                             in_data[88]};
    
    wire lut_731_out = lut_731_table[lut_731_select];
    
    generate
    if ( USE_REG ) begin : ff_731
        reg   lut_731_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_731_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_731_ff <= lut_731_out;
            end
        end
        
        assign out_data[731] = lut_731_ff;
    end
    else begin : no_ff_731
        assign out_data[731] = lut_731_out;
    end
    endgenerate
    
    
    
    // LUT : 732
    wire [63:0] lut_732_table = 64'b0000000000000011000000000000001100000000000000110000000000000011;
    wire [5:0] lut_732_select = {
                             in_data[216],
                             in_data[331],
                             in_data[234],
                             in_data[595],
                             in_data[260],
                             in_data[675]};
    
    wire lut_732_out = lut_732_table[lut_732_select];
    
    generate
    if ( USE_REG ) begin : ff_732
        reg   lut_732_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_732_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_732_ff <= lut_732_out;
            end
        end
        
        assign out_data[732] = lut_732_ff;
    end
    else begin : no_ff_732
        assign out_data[732] = lut_732_out;
    end
    endgenerate
    
    
    
    // LUT : 733
    wire [63:0] lut_733_table = 64'b0010111100001110000010100000100000000100000000000111111101011111;
    wire [5:0] lut_733_select = {
                             in_data[484],
                             in_data[516],
                             in_data[563],
                             in_data[612],
                             in_data[441],
                             in_data[541]};
    
    wire lut_733_out = lut_733_table[lut_733_select];
    
    generate
    if ( USE_REG ) begin : ff_733
        reg   lut_733_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_733_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_733_ff <= lut_733_out;
            end
        end
        
        assign out_data[733] = lut_733_ff;
    end
    else begin : no_ff_733
        assign out_data[733] = lut_733_out;
    end
    endgenerate
    
    
    
    // LUT : 734
    wire [63:0] lut_734_table = 64'b0011001100110011000000000000000000110011001100110000000000000000;
    wire [5:0] lut_734_select = {
                             in_data[692],
                             in_data[497],
                             in_data[460],
                             in_data[363],
                             in_data[683],
                             in_data[724]};
    
    wire lut_734_out = lut_734_table[lut_734_select];
    
    generate
    if ( USE_REG ) begin : ff_734
        reg   lut_734_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_734_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_734_ff <= lut_734_out;
            end
        end
        
        assign out_data[734] = lut_734_ff;
    end
    else begin : no_ff_734
        assign out_data[734] = lut_734_out;
    end
    endgenerate
    
    
    
    // LUT : 735
    wire [63:0] lut_735_table = 64'b1010111111111010101010100000000010101111111111111010101011111010;
    wire [5:0] lut_735_select = {
                             in_data[552],
                             in_data[329],
                             in_data[124],
                             in_data[121],
                             in_data[644],
                             in_data[432]};
    
    wire lut_735_out = lut_735_table[lut_735_select];
    
    generate
    if ( USE_REG ) begin : ff_735
        reg   lut_735_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_735_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_735_ff <= lut_735_out;
            end
        end
        
        assign out_data[735] = lut_735_ff;
    end
    else begin : no_ff_735
        assign out_data[735] = lut_735_out;
    end
    endgenerate
    
    
    
    // LUT : 736
    wire [63:0] lut_736_table = 64'b1100110011001100110011001100110011101110110011001110111011001100;
    wire [5:0] lut_736_select = {
                             in_data[306],
                             in_data[707],
                             in_data[160],
                             in_data[701],
                             in_data[605],
                             in_data[125]};
    
    wire lut_736_out = lut_736_table[lut_736_select];
    
    generate
    if ( USE_REG ) begin : ff_736
        reg   lut_736_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_736_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_736_ff <= lut_736_out;
            end
        end
        
        assign out_data[736] = lut_736_ff;
    end
    else begin : no_ff_736
        assign out_data[736] = lut_736_out;
    end
    endgenerate
    
    
    
    // LUT : 737
    wire [63:0] lut_737_table = 64'b1111111111111111111111111111111111110111001100001111111100110000;
    wire [5:0] lut_737_select = {
                             in_data[249],
                             in_data[561],
                             in_data[492],
                             in_data[401],
                             in_data[382],
                             in_data[67]};
    
    wire lut_737_out = lut_737_table[lut_737_select];
    
    generate
    if ( USE_REG ) begin : ff_737
        reg   lut_737_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_737_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_737_ff <= lut_737_out;
            end
        end
        
        assign out_data[737] = lut_737_ff;
    end
    else begin : no_ff_737
        assign out_data[737] = lut_737_out;
    end
    endgenerate
    
    
    
    // LUT : 738
    wire [63:0] lut_738_table = 64'b1100110011111111000000001011001100000000111111110000000000000000;
    wire [5:0] lut_738_select = {
                             in_data[381],
                             in_data[333],
                             in_data[388],
                             in_data[778],
                             in_data[568],
                             in_data[137]};
    
    wire lut_738_out = lut_738_table[lut_738_select];
    
    generate
    if ( USE_REG ) begin : ff_738
        reg   lut_738_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_738_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_738_ff <= lut_738_out;
            end
        end
        
        assign out_data[738] = lut_738_ff;
    end
    else begin : no_ff_738
        assign out_data[738] = lut_738_out;
    end
    endgenerate
    
    
    
    // LUT : 739
    wire [63:0] lut_739_table = 64'b0000000000000000000000010000000000000000000100010000000100010101;
    wire [5:0] lut_739_select = {
                             in_data[463],
                             in_data[41],
                             in_data[293],
                             in_data[117],
                             in_data[501],
                             in_data[507]};
    
    wire lut_739_out = lut_739_table[lut_739_select];
    
    generate
    if ( USE_REG ) begin : ff_739
        reg   lut_739_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_739_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_739_ff <= lut_739_out;
            end
        end
        
        assign out_data[739] = lut_739_ff;
    end
    else begin : no_ff_739
        assign out_data[739] = lut_739_out;
    end
    endgenerate
    
    
    
    // LUT : 740
    wire [63:0] lut_740_table = 64'b1010000011110000101100001111000011111111111111111111111111111111;
    wire [5:0] lut_740_select = {
                             in_data[465],
                             in_data[309],
                             in_data[89],
                             in_data[633],
                             in_data[335],
                             in_data[263]};
    
    wire lut_740_out = lut_740_table[lut_740_select];
    
    generate
    if ( USE_REG ) begin : ff_740
        reg   lut_740_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_740_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_740_ff <= lut_740_out;
            end
        end
        
        assign out_data[740] = lut_740_ff;
    end
    else begin : no_ff_740
        assign out_data[740] = lut_740_out;
    end
    endgenerate
    
    
    
    // LUT : 741
    wire [63:0] lut_741_table = 64'b0000001011111111000000000011001100100000111111110000000000110011;
    wire [5:0] lut_741_select = {
                             in_data[225],
                             in_data[248],
                             in_data[205],
                             in_data[362],
                             in_data[649],
                             in_data[479]};
    
    wire lut_741_out = lut_741_table[lut_741_select];
    
    generate
    if ( USE_REG ) begin : ff_741
        reg   lut_741_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_741_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_741_ff <= lut_741_out;
            end
        end
        
        assign out_data[741] = lut_741_ff;
    end
    else begin : no_ff_741
        assign out_data[741] = lut_741_out;
    end
    endgenerate
    
    
    
    // LUT : 742
    wire [63:0] lut_742_table = 64'b0000000000000000000000000000000011011111000001011111111101001101;
    wire [5:0] lut_742_select = {
                             in_data[655],
                             in_data[582],
                             in_data[717],
                             in_data[69],
                             in_data[700],
                             in_data[221]};
    
    wire lut_742_out = lut_742_table[lut_742_select];
    
    generate
    if ( USE_REG ) begin : ff_742
        reg   lut_742_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_742_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_742_ff <= lut_742_out;
            end
        end
        
        assign out_data[742] = lut_742_ff;
    end
    else begin : no_ff_742
        assign out_data[742] = lut_742_out;
    end
    endgenerate
    
    
    
    // LUT : 743
    wire [63:0] lut_743_table = 64'b0000111100001111000011110000111100001110000011100000111000001110;
    wire [5:0] lut_743_select = {
                             in_data[386],
                             in_data[32],
                             in_data[45],
                             in_data[93],
                             in_data[742],
                             in_data[262]};
    
    wire lut_743_out = lut_743_table[lut_743_select];
    
    generate
    if ( USE_REG ) begin : ff_743
        reg   lut_743_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_743_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_743_ff <= lut_743_out;
            end
        end
        
        assign out_data[743] = lut_743_ff;
    end
    else begin : no_ff_743
        assign out_data[743] = lut_743_out;
    end
    endgenerate
    
    
    
    // LUT : 744
    wire [63:0] lut_744_table = 64'b0000000011111111000100001111111100000000111111110001000011111111;
    wire [5:0] lut_744_select = {
                             in_data[307],
                             in_data[96],
                             in_data[323],
                             in_data[60],
                             in_data[547],
                             in_data[443]};
    
    wire lut_744_out = lut_744_table[lut_744_select];
    
    generate
    if ( USE_REG ) begin : ff_744
        reg   lut_744_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_744_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_744_ff <= lut_744_out;
            end
        end
        
        assign out_data[744] = lut_744_ff;
    end
    else begin : no_ff_744
        assign out_data[744] = lut_744_out;
    end
    endgenerate
    
    
    
    // LUT : 745
    wire [63:0] lut_745_table = 64'b1010101010101010101010101010101011111111111111111111101011111010;
    wire [5:0] lut_745_select = {
                             in_data[741],
                             in_data[511],
                             in_data[308],
                             in_data[73],
                             in_data[780],
                             in_data[565]};
    
    wire lut_745_out = lut_745_table[lut_745_select];
    
    generate
    if ( USE_REG ) begin : ff_745
        reg   lut_745_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_745_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_745_ff <= lut_745_out;
            end
        end
        
        assign out_data[745] = lut_745_ff;
    end
    else begin : no_ff_745
        assign out_data[745] = lut_745_out;
    end
    endgenerate
    
    
    
    // LUT : 746
    wire [63:0] lut_746_table = 64'b0011001100010011000000000000000010111111101100110000000000000000;
    wire [5:0] lut_746_select = {
                             in_data[546],
                             in_data[487],
                             in_data[614],
                             in_data[251],
                             in_data[192],
                             in_data[592]};
    
    wire lut_746_out = lut_746_table[lut_746_select];
    
    generate
    if ( USE_REG ) begin : ff_746
        reg   lut_746_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_746_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_746_ff <= lut_746_out;
            end
        end
        
        assign out_data[746] = lut_746_ff;
    end
    else begin : no_ff_746
        assign out_data[746] = lut_746_out;
    end
    endgenerate
    
    
    
    // LUT : 747
    wire [63:0] lut_747_table = 64'b1010000010100000101000001010000011111111111111111111111111111111;
    wire [5:0] lut_747_select = {
                             in_data[661],
                             in_data[90],
                             in_data[390],
                             in_data[708],
                             in_data[666],
                             in_data[261]};
    
    wire lut_747_out = lut_747_table[lut_747_select];
    
    generate
    if ( USE_REG ) begin : ff_747
        reg   lut_747_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_747_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_747_ff <= lut_747_out;
            end
        end
        
        assign out_data[747] = lut_747_ff;
    end
    else begin : no_ff_747
        assign out_data[747] = lut_747_out;
    end
    endgenerate
    
    
    
    // LUT : 748
    wire [63:0] lut_748_table = 64'b0101010101110111000100010001000101010101011101110001000100010001;
    wire [5:0] lut_748_select = {
                             in_data[763],
                             in_data[710],
                             in_data[520],
                             in_data[18],
                             in_data[480],
                             in_data[606]};
    
    wire lut_748_out = lut_748_table[lut_748_select];
    
    generate
    if ( USE_REG ) begin : ff_748
        reg   lut_748_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_748_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_748_ff <= lut_748_out;
            end
        end
        
        assign out_data[748] = lut_748_ff;
    end
    else begin : no_ff_748
        assign out_data[748] = lut_748_out;
    end
    endgenerate
    
    
    
    // LUT : 749
    wire [63:0] lut_749_table = 64'b1100110011001100110011011100110011001100110011001100110011001100;
    wire [5:0] lut_749_select = {
                             in_data[715],
                             in_data[376],
                             in_data[631],
                             in_data[781],
                             in_data[328],
                             in_data[684]};
    
    wire lut_749_out = lut_749_table[lut_749_select];
    
    generate
    if ( USE_REG ) begin : ff_749
        reg   lut_749_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_749_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_749_ff <= lut_749_out;
            end
        end
        
        assign out_data[749] = lut_749_ff;
    end
    else begin : no_ff_749
        assign out_data[749] = lut_749_out;
    end
    endgenerate
    
    
    
    // LUT : 750
    wire [63:0] lut_750_table = 64'b1111111111111111111111111111111111111110111111111111000011110000;
    wire [5:0] lut_750_select = {
                             in_data[538],
                             in_data[622],
                             in_data[417],
                             in_data[604],
                             in_data[757],
                             in_data[618]};
    
    wire lut_750_out = lut_750_table[lut_750_select];
    
    generate
    if ( USE_REG ) begin : ff_750
        reg   lut_750_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_750_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_750_ff <= lut_750_out;
            end
        end
        
        assign out_data[750] = lut_750_ff;
    end
    else begin : no_ff_750
        assign out_data[750] = lut_750_out;
    end
    endgenerate
    
    
    
    // LUT : 751
    wire [63:0] lut_751_table = 64'b0000000001010000111111111111100000000000010100001111111111111110;
    wire [5:0] lut_751_select = {
                             in_data[368],
                             in_data[214],
                             in_data[217],
                             in_data[466],
                             in_data[671],
                             in_data[264]};
    
    wire lut_751_out = lut_751_table[lut_751_select];
    
    generate
    if ( USE_REG ) begin : ff_751
        reg   lut_751_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_751_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_751_ff <= lut_751_out;
            end
        end
        
        assign out_data[751] = lut_751_ff;
    end
    else begin : no_ff_751
        assign out_data[751] = lut_751_out;
    end
    endgenerate
    
    
    
    // LUT : 752
    wire [63:0] lut_752_table = 64'b1111110011111100111111101111110011111100111111001111110111111100;
    wire [5:0] lut_752_select = {
                             in_data[782],
                             in_data[759],
                             in_data[681],
                             in_data[345],
                             in_data[508],
                             in_data[391]};
    
    wire lut_752_out = lut_752_table[lut_752_select];
    
    generate
    if ( USE_REG ) begin : ff_752
        reg   lut_752_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_752_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_752_ff <= lut_752_out;
            end
        end
        
        assign out_data[752] = lut_752_ff;
    end
    else begin : no_ff_752
        assign out_data[752] = lut_752_out;
    end
    endgenerate
    
    
    
    // LUT : 753
    wire [63:0] lut_753_table = 64'b0000111000001110111111111111111100001010000010101111111111111111;
    wire [5:0] lut_753_select = {
                             in_data[190],
                             in_data[385],
                             in_data[200],
                             in_data[413],
                             in_data[760],
                             in_data[526]};
    
    wire lut_753_out = lut_753_table[lut_753_select];
    
    generate
    if ( USE_REG ) begin : ff_753
        reg   lut_753_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_753_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_753_ff <= lut_753_out;
            end
        end
        
        assign out_data[753] = lut_753_ff;
    end
    else begin : no_ff_753
        assign out_data[753] = lut_753_out;
    end
    endgenerate
    
    
    
    // LUT : 754
    wire [63:0] lut_754_table = 64'b1111111111111111111111111111111111111111111110101111101111111010;
    wire [5:0] lut_754_select = {
                             in_data[240],
                             in_data[734],
                             in_data[165],
                             in_data[227],
                             in_data[764],
                             in_data[694]};
    
    wire lut_754_out = lut_754_table[lut_754_select];
    
    generate
    if ( USE_REG ) begin : ff_754
        reg   lut_754_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_754_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_754_ff <= lut_754_out;
            end
        end
        
        assign out_data[754] = lut_754_ff;
    end
    else begin : no_ff_754
        assign out_data[754] = lut_754_out;
    end
    endgenerate
    
    
    
    // LUT : 755
    wire [63:0] lut_755_table = 64'b0010101000101010001010100000101000001010000010100000001000000010;
    wire [5:0] lut_755_select = {
                             in_data[56],
                             in_data[674],
                             in_data[532],
                             in_data[471],
                             in_data[75],
                             in_data[374]};
    
    wire lut_755_out = lut_755_table[lut_755_select];
    
    generate
    if ( USE_REG ) begin : ff_755
        reg   lut_755_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_755_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_755_ff <= lut_755_out;
            end
        end
        
        assign out_data[755] = lut_755_ff;
    end
    else begin : no_ff_755
        assign out_data[755] = lut_755_out;
    end
    endgenerate
    
    
    
    // LUT : 756
    wire [63:0] lut_756_table = 64'b0000000000000000000000000001010100000000000000000000000000010101;
    wire [5:0] lut_756_select = {
                             in_data[337],
                             in_data[464],
                             in_data[743],
                             in_data[313],
                             in_data[726],
                             in_data[294]};
    
    wire lut_756_out = lut_756_table[lut_756_select];
    
    generate
    if ( USE_REG ) begin : ff_756
        reg   lut_756_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_756_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_756_ff <= lut_756_out;
            end
        end
        
        assign out_data[756] = lut_756_ff;
    end
    else begin : no_ff_756
        assign out_data[756] = lut_756_out;
    end
    endgenerate
    
    
    
    // LUT : 757
    wire [63:0] lut_757_table = 64'b1100110011001100111011101111111011001100110011001110111011101110;
    wire [5:0] lut_757_select = {
                             in_data[779],
                             in_data[722],
                             in_data[61],
                             in_data[7],
                             in_data[593],
                             in_data[230]};
    
    wire lut_757_out = lut_757_table[lut_757_select];
    
    generate
    if ( USE_REG ) begin : ff_757
        reg   lut_757_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_757_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_757_ff <= lut_757_out;
            end
        end
        
        assign out_data[757] = lut_757_ff;
    end
    else begin : no_ff_757
        assign out_data[757] = lut_757_out;
    end
    endgenerate
    
    
    
    // LUT : 758
    wire [63:0] lut_758_table = 64'b1111111111111111111111111111111111111111111111111010101010101010;
    wire [5:0] lut_758_select = {
                             in_data[680],
                             in_data[370],
                             in_data[84],
                             in_data[698],
                             in_data[616],
                             in_data[167]};
    
    wire lut_758_out = lut_758_table[lut_758_select];
    
    generate
    if ( USE_REG ) begin : ff_758
        reg   lut_758_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_758_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_758_ff <= lut_758_out;
            end
        end
        
        assign out_data[758] = lut_758_ff;
    end
    else begin : no_ff_758
        assign out_data[758] = lut_758_out;
    end
    endgenerate
    
    
    
    // LUT : 759
    wire [63:0] lut_759_table = 64'b1111110011111100110111001101110011111100111111001101110011011100;
    wire [5:0] lut_759_select = {
                             in_data[736],
                             in_data[177],
                             in_data[116],
                             in_data[322],
                             in_data[677],
                             in_data[657]};
    
    wire lut_759_out = lut_759_table[lut_759_select];
    
    generate
    if ( USE_REG ) begin : ff_759
        reg   lut_759_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_759_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_759_ff <= lut_759_out;
            end
        end
        
        assign out_data[759] = lut_759_ff;
    end
    else begin : no_ff_759
        assign out_data[759] = lut_759_out;
    end
    endgenerate
    
    
    
    // LUT : 760
    wire [63:0] lut_760_table = 64'b0000000000000000000000000111111100000000000011110000111101111111;
    wire [5:0] lut_760_select = {
                             in_data[650],
                             in_data[274],
                             in_data[349],
                             in_data[318],
                             in_data[758],
                             in_data[166]};
    
    wire lut_760_out = lut_760_table[lut_760_select];
    
    generate
    if ( USE_REG ) begin : ff_760
        reg   lut_760_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_760_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_760_ff <= lut_760_out;
            end
        end
        
        assign out_data[760] = lut_760_ff;
    end
    else begin : no_ff_760
        assign out_data[760] = lut_760_out;
    end
    endgenerate
    
    
    
    // LUT : 761
    wire [63:0] lut_761_table = 64'b0000001010101011000000000010101100000000001010110000000000101011;
    wire [5:0] lut_761_select = {
                             in_data[62],
                             in_data[783],
                             in_data[549],
                             in_data[127],
                             in_data[474],
                             in_data[705]};
    
    wire lut_761_out = lut_761_table[lut_761_select];
    
    generate
    if ( USE_REG ) begin : ff_761
        reg   lut_761_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_761_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_761_ff <= lut_761_out;
            end
        end
        
        assign out_data[761] = lut_761_ff;
    end
    else begin : no_ff_761
        assign out_data[761] = lut_761_out;
    end
    endgenerate
    
    
    
    // LUT : 762
    wire [63:0] lut_762_table = 64'b1111111111111111111111111111111110101010101010101010101010101010;
    wire [5:0] lut_762_select = {
                             in_data[713],
                             in_data[718],
                             in_data[6],
                             in_data[344],
                             in_data[395],
                             in_data[553]};
    
    wire lut_762_out = lut_762_table[lut_762_select];
    
    generate
    if ( USE_REG ) begin : ff_762
        reg   lut_762_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_762_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_762_ff <= lut_762_out;
            end
        end
        
        assign out_data[762] = lut_762_ff;
    end
    else begin : no_ff_762
        assign out_data[762] = lut_762_out;
    end
    endgenerate
    
    
    
    // LUT : 763
    wire [63:0] lut_763_table = 64'b1111111111111111111111101111101011111111111100101111111011110010;
    wire [5:0] lut_763_select = {
                             in_data[371],
                             in_data[91],
                             in_data[427],
                             in_data[100],
                             in_data[191],
                             in_data[433]};
    
    wire lut_763_out = lut_763_table[lut_763_select];
    
    generate
    if ( USE_REG ) begin : ff_763
        reg   lut_763_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_763_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_763_ff <= lut_763_out;
            end
        end
        
        assign out_data[763] = lut_763_ff;
    end
    else begin : no_ff_763
        assign out_data[763] = lut_763_out;
    end
    endgenerate
    
    
    
    // LUT : 764
    wire [63:0] lut_764_table = 64'b0101110100000000111111111010101011010101000000001111111110101010;
    wire [5:0] lut_764_select = {
                             in_data[278],
                             in_data[404],
                             in_data[523],
                             in_data[531],
                             in_data[28],
                             in_data[146]};
    
    wire lut_764_out = lut_764_table[lut_764_select];
    
    generate
    if ( USE_REG ) begin : ff_764
        reg   lut_764_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_764_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_764_ff <= lut_764_out;
            end
        end
        
        assign out_data[764] = lut_764_ff;
    end
    else begin : no_ff_764
        assign out_data[764] = lut_764_out;
    end
    endgenerate
    
    
    
    // LUT : 765
    wire [63:0] lut_765_table = 64'b0000000000001111000000000000000000001111111111110000000000001111;
    wire [5:0] lut_765_select = {
                             in_data[745],
                             in_data[129],
                             in_data[744],
                             in_data[235],
                             in_data[560],
                             in_data[559]};
    
    wire lut_765_out = lut_765_table[lut_765_select];
    
    generate
    if ( USE_REG ) begin : ff_765
        reg   lut_765_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_765_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_765_ff <= lut_765_out;
            end
        end
        
        assign out_data[765] = lut_765_ff;
    end
    else begin : no_ff_765
        assign out_data[765] = lut_765_out;
    end
    endgenerate
    
    
    
    // LUT : 766
    wire [63:0] lut_766_table = 64'b1100110011001100111111111111111100000100000001001100110111001101;
    wire [5:0] lut_766_select = {
                             in_data[277],
                             in_data[534],
                             in_data[725],
                             in_data[178],
                             in_data[193],
                             in_data[586]};
    
    wire lut_766_out = lut_766_table[lut_766_select];
    
    generate
    if ( USE_REG ) begin : ff_766
        reg   lut_766_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_766_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_766_ff <= lut_766_out;
            end
        end
        
        assign out_data[766] = lut_766_ff;
    end
    else begin : no_ff_766
        assign out_data[766] = lut_766_out;
    end
    endgenerate
    
    
    
    // LUT : 767
    wire [63:0] lut_767_table = 64'b0000111100001111000011000000110000001111000011110000110000001100;
    wire [5:0] lut_767_select = {
                             in_data[754],
                             in_data[312],
                             in_data[48],
                             in_data[749],
                             in_data[194],
                             in_data[420]};
    
    wire lut_767_out = lut_767_table[lut_767_select];
    
    generate
    if ( USE_REG ) begin : ff_767
        reg   lut_767_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_767_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_767_ff <= lut_767_out;
            end
        end
        
        assign out_data[767] = lut_767_ff;
    end
    else begin : no_ff_767
        assign out_data[767] = lut_767_out;
    end
    endgenerate
    
    
    
    // LUT : 768
    wire [63:0] lut_768_table = 64'b1101010111010101010001010100010111000101110001010100010101000101;
    wire [5:0] lut_768_select = {
                             in_data[222],
                             in_data[279],
                             in_data[34],
                             in_data[435],
                             in_data[285],
                             in_data[131]};
    
    wire lut_768_out = lut_768_table[lut_768_select];
    
    generate
    if ( USE_REG ) begin : ff_768
        reg   lut_768_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_768_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_768_ff <= lut_768_out;
            end
        end
        
        assign out_data[768] = lut_768_ff;
    end
    else begin : no_ff_768
        assign out_data[768] = lut_768_out;
    end
    endgenerate
    
    
    
    // LUT : 769
    wire [63:0] lut_769_table = 64'b1100110011001100111011101110110011001100110011001110110011111100;
    wire [5:0] lut_769_select = {
                             in_data[336],
                             in_data[408],
                             in_data[55],
                             in_data[639],
                             in_data[350],
                             in_data[591]};
    
    wire lut_769_out = lut_769_table[lut_769_select];
    
    generate
    if ( USE_REG ) begin : ff_769
        reg   lut_769_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_769_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_769_ff <= lut_769_out;
            end
        end
        
        assign out_data[769] = lut_769_ff;
    end
    else begin : no_ff_769
        assign out_data[769] = lut_769_out;
    end
    endgenerate
    
    
    
    // LUT : 770
    wire [63:0] lut_770_table = 64'b0111011101110111001100110011001100110001001100000011000100110000;
    wire [5:0] lut_770_select = {
                             in_data[346],
                             in_data[184],
                             in_data[558],
                             in_data[714],
                             in_data[297],
                             in_data[321]};
    
    wire lut_770_out = lut_770_table[lut_770_select];
    
    generate
    if ( USE_REG ) begin : ff_770
        reg   lut_770_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_770_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_770_ff <= lut_770_out;
            end
        end
        
        assign out_data[770] = lut_770_ff;
    end
    else begin : no_ff_770
        assign out_data[770] = lut_770_out;
    end
    endgenerate
    
    
    
    // LUT : 771
    wire [63:0] lut_771_table = 64'b1111111111111111111111111111111111111110111111001111111011111100;
    wire [5:0] lut_771_select = {
                             in_data[66],
                             in_data[81],
                             in_data[25],
                             in_data[416],
                             in_data[607],
                             in_data[280]};
    
    wire lut_771_out = lut_771_table[lut_771_select];
    
    generate
    if ( USE_REG ) begin : ff_771
        reg   lut_771_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_771_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_771_ff <= lut_771_out;
            end
        end
        
        assign out_data[771] = lut_771_ff;
    end
    else begin : no_ff_771
        assign out_data[771] = lut_771_out;
    end
    endgenerate
    
    
    
    // LUT : 772
    wire [63:0] lut_772_table = 64'b1010000010101010001000101010101000000000111110100010001011111111;
    wire [5:0] lut_772_select = {
                             in_data[245],
                             in_data[197],
                             in_data[304],
                             in_data[421],
                             in_data[762],
                             in_data[103]};
    
    wire lut_772_out = lut_772_table[lut_772_select];
    
    generate
    if ( USE_REG ) begin : ff_772
        reg   lut_772_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_772_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_772_ff <= lut_772_out;
            end
        end
        
        assign out_data[772] = lut_772_ff;
    end
    else begin : no_ff_772
        assign out_data[772] = lut_772_out;
    end
    endgenerate
    
    
    
    // LUT : 773
    wire [63:0] lut_773_table = 64'b0100110000000000000000000000000011111111010101011101110101010101;
    wire [5:0] lut_773_select = {
                             in_data[536],
                             in_data[78],
                             in_data[665],
                             in_data[86],
                             in_data[288],
                             in_data[498]};
    
    wire lut_773_out = lut_773_table[lut_773_select];
    
    generate
    if ( USE_REG ) begin : ff_773
        reg   lut_773_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_773_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_773_ff <= lut_773_out;
            end
        end
        
        assign out_data[773] = lut_773_ff;
    end
    else begin : no_ff_773
        assign out_data[773] = lut_773_out;
    end
    endgenerate
    
    
    
    // LUT : 774
    wire [63:0] lut_774_table = 64'b0000000000001110000001000000111110000100100011101000110011001110;
    wire [5:0] lut_774_select = {
                             in_data[429],
                             in_data[678],
                             in_data[272],
                             in_data[298],
                             in_data[237],
                             in_data[290]};
    
    wire lut_774_out = lut_774_table[lut_774_select];
    
    generate
    if ( USE_REG ) begin : ff_774
        reg   lut_774_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_774_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_774_ff <= lut_774_out;
            end
        end
        
        assign out_data[774] = lut_774_ff;
    end
    else begin : no_ff_774
        assign out_data[774] = lut_774_out;
    end
    endgenerate
    
    
    
    // LUT : 775
    wire [63:0] lut_775_table = 64'b1111000011110000111111111111010110100000101000001111111111111111;
    wire [5:0] lut_775_select = {
                             in_data[510],
                             in_data[210],
                             in_data[777],
                             in_data[172],
                             in_data[198],
                             in_data[621]};
    
    wire lut_775_out = lut_775_table[lut_775_select];
    
    generate
    if ( USE_REG ) begin : ff_775
        reg   lut_775_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_775_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_775_ff <= lut_775_out;
            end
        end
        
        assign out_data[775] = lut_775_ff;
    end
    else begin : no_ff_775
        assign out_data[775] = lut_775_out;
    end
    endgenerate
    
    
    
    // LUT : 776
    wire [63:0] lut_776_table = 64'b1100110000000000111111111100000011001100000000001111111111001000;
    wire [5:0] lut_776_select = {
                             in_data[447],
                             in_data[446],
                             in_data[470],
                             in_data[765],
                             in_data[373],
                             in_data[195]};
    
    wire lut_776_out = lut_776_table[lut_776_select];
    
    generate
    if ( USE_REG ) begin : ff_776
        reg   lut_776_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_776_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_776_ff <= lut_776_out;
            end
        end
        
        assign out_data[776] = lut_776_ff;
    end
    else begin : no_ff_776
        assign out_data[776] = lut_776_out;
    end
    endgenerate
    
    
    
    // LUT : 777
    wire [63:0] lut_777_table = 64'b1101000011000000111111011111110011010100110000001111111111111101;
    wire [5:0] lut_777_select = {
                             in_data[188],
                             in_data[295],
                             in_data[693],
                             in_data[467],
                             in_data[163],
                             in_data[690]};
    
    wire lut_777_out = lut_777_table[lut_777_select];
    
    generate
    if ( USE_REG ) begin : ff_777
        reg   lut_777_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_777_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_777_ff <= lut_777_out;
            end
        end
        
        assign out_data[777] = lut_777_ff;
    end
    else begin : no_ff_777
        assign out_data[777] = lut_777_out;
    end
    endgenerate
    
    
    
    // LUT : 778
    wire [63:0] lut_778_table = 64'b1111110011111100111111001111111111111100111111001111111011111100;
    wire [5:0] lut_778_select = {
                             in_data[1],
                             in_data[327],
                             in_data[751],
                             in_data[130],
                             in_data[554],
                             in_data[283]};
    
    wire lut_778_out = lut_778_table[lut_778_select];
    
    generate
    if ( USE_REG ) begin : ff_778
        reg   lut_778_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_778_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_778_ff <= lut_778_out;
            end
        end
        
        assign out_data[778] = lut_778_ff;
    end
    else begin : no_ff_778
        assign out_data[778] = lut_778_out;
    end
    endgenerate
    
    
    
    // LUT : 779
    wire [63:0] lut_779_table = 64'b1110000010000000111110001111111111100000101000001111101011111111;
    wire [5:0] lut_779_select = {
                             in_data[449],
                             in_data[496],
                             in_data[454],
                             in_data[584],
                             in_data[589],
                             in_data[585]};
    
    wire lut_779_out = lut_779_table[lut_779_select];
    
    generate
    if ( USE_REG ) begin : ff_779
        reg   lut_779_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_779_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_779_ff <= lut_779_out;
            end
        end
        
        assign out_data[779] = lut_779_ff;
    end
    else begin : no_ff_779
        assign out_data[779] = lut_779_out;
    end
    endgenerate
    
    
    
    // LUT : 780
    wire [63:0] lut_780_table = 64'b0000001100000001111111111111010011111111111100111111110001110100;
    wire [5:0] lut_780_select = {
                             in_data[509],
                             in_data[551],
                             in_data[361],
                             in_data[571],
                             in_data[300],
                             in_data[620]};
    
    wire lut_780_out = lut_780_table[lut_780_select];
    
    generate
    if ( USE_REG ) begin : ff_780
        reg   lut_780_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_780_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_780_ff <= lut_780_out;
            end
        end
        
        assign out_data[780] = lut_780_ff;
    end
    else begin : no_ff_780
        assign out_data[780] = lut_780_out;
    end
    endgenerate
    
    
    
    // LUT : 781
    wire [63:0] lut_781_table = 64'b0000110000001111000000000000111100001100000011110000000000001111;
    wire [5:0] lut_781_select = {
                             in_data[756],
                             in_data[697],
                             in_data[449],
                             in_data[397],
                             in_data[170],
                             in_data[33]};
    
    wire lut_781_out = lut_781_table[lut_781_select];
    
    generate
    if ( USE_REG ) begin : ff_781
        reg   lut_781_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_781_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_781_ff <= lut_781_out;
            end
        end
        
        assign out_data[781] = lut_781_ff;
    end
    else begin : no_ff_781
        assign out_data[781] = lut_781_out;
    end
    endgenerate
    
    
    
    // LUT : 782
    wire [63:0] lut_782_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_782_select = {
                             in_data[485],
                             in_data[194],
                             in_data[184],
                             in_data[562],
                             in_data[779],
                             in_data[614]};
    
    wire lut_782_out = lut_782_table[lut_782_select];
    
    generate
    if ( USE_REG ) begin : ff_782
        reg   lut_782_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_782_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_782_ff <= lut_782_out;
            end
        end
        
        assign out_data[782] = lut_782_ff;
    end
    else begin : no_ff_782
        assign out_data[782] = lut_782_out;
    end
    endgenerate
    
    
    
    // LUT : 783
    wire [63:0] lut_783_table = 64'b0000000000000000010101010101000111010101110101011111111111111111;
    wire [5:0] lut_783_select = {
                             in_data[352],
                             in_data[427],
                             in_data[111],
                             in_data[603],
                             in_data[52],
                             in_data[215]};
    
    wire lut_783_out = lut_783_table[lut_783_select];
    
    generate
    if ( USE_REG ) begin : ff_783
        reg   lut_783_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_783_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_783_ff <= lut_783_out;
            end
        end
        
        assign out_data[783] = lut_783_ff;
    end
    else begin : no_ff_783
        assign out_data[783] = lut_783_out;
    end
    endgenerate
    
    
    
    // LUT : 784
    wire [63:0] lut_784_table = 64'b0000000011101110000000000000000001010101111101010101010101010101;
    wire [5:0] lut_784_select = {
                             in_data[434],
                             in_data[520],
                             in_data[557],
                             in_data[76],
                             in_data[506],
                             in_data[403]};
    
    wire lut_784_out = lut_784_table[lut_784_select];
    
    generate
    if ( USE_REG ) begin : ff_784
        reg   lut_784_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_784_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_784_ff <= lut_784_out;
            end
        end
        
        assign out_data[784] = lut_784_ff;
    end
    else begin : no_ff_784
        assign out_data[784] = lut_784_out;
    end
    endgenerate
    
    
    
    // LUT : 785
    wire [63:0] lut_785_table = 64'b0001000100110010001100111011101100010001001000000011001110111011;
    wire [5:0] lut_785_select = {
                             in_data[418],
                             in_data[425],
                             in_data[469],
                             in_data[761],
                             in_data[213],
                             in_data[541]};
    
    wire lut_785_out = lut_785_table[lut_785_select];
    
    generate
    if ( USE_REG ) begin : ff_785
        reg   lut_785_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_785_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_785_ff <= lut_785_out;
            end
        end
        
        assign out_data[785] = lut_785_ff;
    end
    else begin : no_ff_785
        assign out_data[785] = lut_785_out;
    end
    endgenerate
    
    
    
    // LUT : 786
    wire [63:0] lut_786_table = 64'b0000000000000000001100110011001100000000000000000011000000110011;
    wire [5:0] lut_786_select = {
                             in_data[676],
                             in_data[190],
                             in_data[71],
                             in_data[438],
                             in_data[130],
                             in_data[753]};
    
    wire lut_786_out = lut_786_table[lut_786_select];
    
    generate
    if ( USE_REG ) begin : ff_786
        reg   lut_786_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_786_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_786_ff <= lut_786_out;
            end
        end
        
        assign out_data[786] = lut_786_ff;
    end
    else begin : no_ff_786
        assign out_data[786] = lut_786_out;
    end
    endgenerate
    
    
    
    // LUT : 787
    wire [63:0] lut_787_table = 64'b1111010111110101010100010101000111110101111101010101000001010001;
    wire [5:0] lut_787_select = {
                             in_data[226],
                             in_data[273],
                             in_data[759],
                             in_data[341],
                             in_data[724],
                             in_data[159]};
    
    wire lut_787_out = lut_787_table[lut_787_select];
    
    generate
    if ( USE_REG ) begin : ff_787
        reg   lut_787_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_787_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_787_ff <= lut_787_out;
            end
        end
        
        assign out_data[787] = lut_787_ff;
    end
    else begin : no_ff_787
        assign out_data[787] = lut_787_out;
    end
    endgenerate
    
    
    
    // LUT : 788
    wire [63:0] lut_788_table = 64'b0010111000000111101011100000111111111111000000001111111100000000;
    wire [5:0] lut_788_select = {
                             in_data[483],
                             in_data[54],
                             in_data[486],
                             in_data[678],
                             in_data[390],
                             in_data[85]};
    
    wire lut_788_out = lut_788_table[lut_788_select];
    
    generate
    if ( USE_REG ) begin : ff_788
        reg   lut_788_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_788_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_788_ff <= lut_788_out;
            end
        end
        
        assign out_data[788] = lut_788_ff;
    end
    else begin : no_ff_788
        assign out_data[788] = lut_788_out;
    end
    endgenerate
    
    
    
    // LUT : 789
    wire [63:0] lut_789_table = 64'b0101011100000000010111110101011100010001000000000101010100000001;
    wire [5:0] lut_789_select = {
                             in_data[655],
                             in_data[460],
                             in_data[208],
                             in_data[380],
                             in_data[635],
                             in_data[578]};
    
    wire lut_789_out = lut_789_table[lut_789_select];
    
    generate
    if ( USE_REG ) begin : ff_789
        reg   lut_789_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_789_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_789_ff <= lut_789_out;
            end
        end
        
        assign out_data[789] = lut_789_ff;
    end
    else begin : no_ff_789
        assign out_data[789] = lut_789_out;
    end
    endgenerate
    
    
    
    // LUT : 790
    wire [63:0] lut_790_table = 64'b1100111011011110100011111100111111111110111111101100111111001111;
    wire [5:0] lut_790_select = {
                             in_data[14],
                             in_data[294],
                             in_data[223],
                             in_data[349],
                             in_data[712],
                             in_data[684]};
    
    wire lut_790_out = lut_790_table[lut_790_select];
    
    generate
    if ( USE_REG ) begin : ff_790
        reg   lut_790_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_790_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_790_ff <= lut_790_out;
            end
        end
        
        assign out_data[790] = lut_790_ff;
    end
    else begin : no_ff_790
        assign out_data[790] = lut_790_out;
    end
    endgenerate
    
    
    
    // LUT : 791
    wire [63:0] lut_791_table = 64'b1010101000000000111011101000100011111111111011101111111111101110;
    wire [5:0] lut_791_select = {
                             in_data[720],
                             in_data[140],
                             in_data[677],
                             in_data[27],
                             in_data[394],
                             in_data[735]};
    
    wire lut_791_out = lut_791_table[lut_791_select];
    
    generate
    if ( USE_REG ) begin : ff_791
        reg   lut_791_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_791_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_791_ff <= lut_791_out;
            end
        end
        
        assign out_data[791] = lut_791_ff;
    end
    else begin : no_ff_791
        assign out_data[791] = lut_791_out;
    end
    endgenerate
    
    
    
    // LUT : 792
    wire [63:0] lut_792_table = 64'b1110111011111111111011111111111111001110111011111100111011101110;
    wire [5:0] lut_792_select = {
                             in_data[563],
                             in_data[758],
                             in_data[286],
                             in_data[502],
                             in_data[387],
                             in_data[276]};
    
    wire lut_792_out = lut_792_table[lut_792_select];
    
    generate
    if ( USE_REG ) begin : ff_792
        reg   lut_792_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_792_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_792_ff <= lut_792_out;
            end
        end
        
        assign out_data[792] = lut_792_ff;
    end
    else begin : no_ff_792
        assign out_data[792] = lut_792_out;
    end
    endgenerate
    
    
    
    // LUT : 793
    wire [63:0] lut_793_table = 64'b1111111111111111111111110000111111111111111111111101111100001111;
    wire [5:0] lut_793_select = {
                             in_data[499],
                             in_data[135],
                             in_data[611],
                             in_data[428],
                             in_data[302],
                             in_data[778]};
    
    wire lut_793_out = lut_793_table[lut_793_select];
    
    generate
    if ( USE_REG ) begin : ff_793
        reg   lut_793_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_793_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_793_ff <= lut_793_out;
            end
        end
        
        assign out_data[793] = lut_793_ff;
    end
    else begin : no_ff_793
        assign out_data[793] = lut_793_out;
    end
    endgenerate
    
    
    
    // LUT : 794
    wire [63:0] lut_794_table = 64'b0001110111011101000100010001100101011101100110010001100100011001;
    wire [5:0] lut_794_select = {
                             in_data[24],
                             in_data[311],
                             in_data[112],
                             in_data[391],
                             in_data[429],
                             in_data[455]};
    
    wire lut_794_out = lut_794_table[lut_794_select];
    
    generate
    if ( USE_REG ) begin : ff_794
        reg   lut_794_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_794_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_794_ff <= lut_794_out;
            end
        end
        
        assign out_data[794] = lut_794_ff;
    end
    else begin : no_ff_794
        assign out_data[794] = lut_794_out;
    end
    endgenerate
    
    
    
    // LUT : 795
    wire [63:0] lut_795_table = 64'b1111001111110011111100101111001011110011111100111111001011110010;
    wire [5:0] lut_795_select = {
                             in_data[30],
                             in_data[439],
                             in_data[84],
                             in_data[480],
                             in_data[315],
                             in_data[13]};
    
    wire lut_795_out = lut_795_table[lut_795_select];
    
    generate
    if ( USE_REG ) begin : ff_795
        reg   lut_795_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_795_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_795_ff <= lut_795_out;
            end
        end
        
        assign out_data[795] = lut_795_ff;
    end
    else begin : no_ff_795
        assign out_data[795] = lut_795_out;
    end
    endgenerate
    
    
    
    // LUT : 796
    wire [63:0] lut_796_table = 64'b0000000001010101000000000101010100000000000100000000000001010101;
    wire [5:0] lut_796_select = {
                             in_data[309],
                             in_data[612],
                             in_data[229],
                             in_data[703],
                             in_data[437],
                             in_data[123]};
    
    wire lut_796_out = lut_796_table[lut_796_select];
    
    generate
    if ( USE_REG ) begin : ff_796
        reg   lut_796_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_796_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_796_ff <= lut_796_out;
            end
        end
        
        assign out_data[796] = lut_796_ff;
    end
    else begin : no_ff_796
        assign out_data[796] = lut_796_out;
    end
    endgenerate
    
    
    
    // LUT : 797
    wire [63:0] lut_797_table = 64'b1111111111111110111111111111111111111111111111101111111011111110;
    wire [5:0] lut_797_select = {
                             in_data[269],
                             in_data[161],
                             in_data[743],
                             in_data[136],
                             in_data[535],
                             in_data[651]};
    
    wire lut_797_out = lut_797_table[lut_797_select];
    
    generate
    if ( USE_REG ) begin : ff_797
        reg   lut_797_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_797_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_797_ff <= lut_797_out;
            end
        end
        
        assign out_data[797] = lut_797_ff;
    end
    else begin : no_ff_797
        assign out_data[797] = lut_797_out;
    end
    endgenerate
    
    
    
    // LUT : 798
    wire [63:0] lut_798_table = 64'b1111101011111111111110001111111100000000010101000000000001010101;
    wire [5:0] lut_798_select = {
                             in_data[266],
                             in_data[306],
                             in_data[262],
                             in_data[322],
                             in_data[285],
                             in_data[316]};
    
    wire lut_798_out = lut_798_table[lut_798_select];
    
    generate
    if ( USE_REG ) begin : ff_798
        reg   lut_798_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_798_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_798_ff <= lut_798_out;
            end
        end
        
        assign out_data[798] = lut_798_ff;
    end
    else begin : no_ff_798
        assign out_data[798] = lut_798_out;
    end
    endgenerate
    
    
    
    // LUT : 799
    wire [63:0] lut_799_table = 64'b1111000000100000111100001111000011110000111100001111000011111010;
    wire [5:0] lut_799_select = {
                             in_data[171],
                             in_data[228],
                             in_data[622],
                             in_data[128],
                             in_data[141],
                             in_data[443]};
    
    wire lut_799_out = lut_799_table[lut_799_select];
    
    generate
    if ( USE_REG ) begin : ff_799
        reg   lut_799_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_799_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_799_ff <= lut_799_out;
            end
        end
        
        assign out_data[799] = lut_799_ff;
    end
    else begin : no_ff_799
        assign out_data[799] = lut_799_out;
    end
    endgenerate
    
    
    
    // LUT : 800
    wire [63:0] lut_800_table = 64'b0000111100001111000000110000111100001111000011110000001100001111;
    wire [5:0] lut_800_select = {
                             in_data[82],
                             in_data[156],
                             in_data[771],
                             in_data[290],
                             in_data[3],
                             in_data[644]};
    
    wire lut_800_out = lut_800_table[lut_800_select];
    
    generate
    if ( USE_REG ) begin : ff_800
        reg   lut_800_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_800_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_800_ff <= lut_800_out;
            end
        end
        
        assign out_data[800] = lut_800_ff;
    end
    else begin : no_ff_800
        assign out_data[800] = lut_800_out;
    end
    endgenerate
    
    
    
    // LUT : 801
    wire [63:0] lut_801_table = 64'b0000000000000000000000000000000000000001010011110000000001001111;
    wire [5:0] lut_801_select = {
                             in_data[625],
                             in_data[531],
                             in_data[683],
                             in_data[544],
                             in_data[230],
                             in_data[92]};
    
    wire lut_801_out = lut_801_table[lut_801_select];
    
    generate
    if ( USE_REG ) begin : ff_801
        reg   lut_801_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_801_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_801_ff <= lut_801_out;
            end
        end
        
        assign out_data[801] = lut_801_ff;
    end
    else begin : no_ff_801
        assign out_data[801] = lut_801_out;
    end
    endgenerate
    
    
    
    // LUT : 802
    wire [63:0] lut_802_table = 64'b0000100011101110000000000000000010001000111011100000000011001100;
    wire [5:0] lut_802_select = {
                             in_data[479],
                             in_data[324],
                             in_data[685],
                             in_data[166],
                             in_data[410],
                             in_data[621]};
    
    wire lut_802_out = lut_802_table[lut_802_select];
    
    generate
    if ( USE_REG ) begin : ff_802
        reg   lut_802_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_802_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_802_ff <= lut_802_out;
            end
        end
        
        assign out_data[802] = lut_802_ff;
    end
    else begin : no_ff_802
        assign out_data[802] = lut_802_out;
    end
    endgenerate
    
    
    
    // LUT : 803
    wire [63:0] lut_803_table = 64'b1111111111111111111111111111111111101110111011101110111011101110;
    wire [5:0] lut_803_select = {
                             in_data[649],
                             in_data[670],
                             in_data[601],
                             in_data[250],
                             in_data[664],
                             in_data[323]};
    
    wire lut_803_out = lut_803_table[lut_803_select];
    
    generate
    if ( USE_REG ) begin : ff_803
        reg   lut_803_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_803_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_803_ff <= lut_803_out;
            end
        end
        
        assign out_data[803] = lut_803_ff;
    end
    else begin : no_ff_803
        assign out_data[803] = lut_803_out;
    end
    endgenerate
    
    
    
    // LUT : 804
    wire [63:0] lut_804_table = 64'b1100110011001100110011001110111011001110111011101000100010001000;
    wire [5:0] lut_804_select = {
                             in_data[371],
                             in_data[291],
                             in_data[476],
                             in_data[86],
                             in_data[546],
                             in_data[426]};
    
    wire lut_804_out = lut_804_table[lut_804_select];
    
    generate
    if ( USE_REG ) begin : ff_804
        reg   lut_804_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_804_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_804_ff <= lut_804_out;
            end
        end
        
        assign out_data[804] = lut_804_ff;
    end
    else begin : no_ff_804
        assign out_data[804] = lut_804_out;
    end
    endgenerate
    
    
    
    // LUT : 805
    wire [63:0] lut_805_table = 64'b0101000100010001000100010001001100000000001000000000000000000000;
    wire [5:0] lut_805_select = {
                             in_data[490],
                             in_data[67],
                             in_data[16],
                             in_data[393],
                             in_data[717],
                             in_data[628]};
    
    wire lut_805_out = lut_805_table[lut_805_select];
    
    generate
    if ( USE_REG ) begin : ff_805
        reg   lut_805_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_805_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_805_ff <= lut_805_out;
            end
        end
        
        assign out_data[805] = lut_805_ff;
    end
    else begin : no_ff_805
        assign out_data[805] = lut_805_out;
    end
    endgenerate
    
    
    
    // LUT : 806
    wire [63:0] lut_806_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_806_select = {
                             in_data[210],
                             in_data[53],
                             in_data[591],
                             in_data[8],
                             in_data[671],
                             in_data[150]};
    
    wire lut_806_out = lut_806_table[lut_806_select];
    
    generate
    if ( USE_REG ) begin : ff_806
        reg   lut_806_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_806_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_806_ff <= lut_806_out;
            end
        end
        
        assign out_data[806] = lut_806_ff;
    end
    else begin : no_ff_806
        assign out_data[806] = lut_806_out;
    end
    endgenerate
    
    
    
    // LUT : 807
    wire [63:0] lut_807_table = 64'b1111111111110001111100001111000011111111111100111011000011110000;
    wire [5:0] lut_807_select = {
                             in_data[217],
                             in_data[408],
                             in_data[414],
                             in_data[398],
                             in_data[244],
                             in_data[451]};
    
    wire lut_807_out = lut_807_table[lut_807_select];
    
    generate
    if ( USE_REG ) begin : ff_807
        reg   lut_807_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_807_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_807_ff <= lut_807_out;
            end
        end
        
        assign out_data[807] = lut_807_ff;
    end
    else begin : no_ff_807
        assign out_data[807] = lut_807_out;
    end
    endgenerate
    
    
    
    // LUT : 808
    wire [63:0] lut_808_table = 64'b0010001000100010000000000000000011101111001110110000000011111111;
    wire [5:0] lut_808_select = {
                             in_data[180],
                             in_data[293],
                             in_data[234],
                             in_data[584],
                             in_data[399],
                             in_data[609]};
    
    wire lut_808_out = lut_808_table[lut_808_select];
    
    generate
    if ( USE_REG ) begin : ff_808
        reg   lut_808_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_808_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_808_ff <= lut_808_out;
            end
        end
        
        assign out_data[808] = lut_808_ff;
    end
    else begin : no_ff_808
        assign out_data[808] = lut_808_out;
    end
    endgenerate
    
    
    
    // LUT : 809
    wire [63:0] lut_809_table = 64'b1111111111111110111111111111111111111111111111101111111111111110;
    wire [5:0] lut_809_select = {
                             in_data[705],
                             in_data[627],
                             in_data[608],
                             in_data[218],
                             in_data[507],
                             in_data[219]};
    
    wire lut_809_out = lut_809_table[lut_809_select];
    
    generate
    if ( USE_REG ) begin : ff_809
        reg   lut_809_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_809_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_809_ff <= lut_809_out;
            end
        end
        
        assign out_data[809] = lut_809_ff;
    end
    else begin : no_ff_809
        assign out_data[809] = lut_809_out;
    end
    endgenerate
    
    
    
    // LUT : 810
    wire [63:0] lut_810_table = 64'b1111111111101100111111111111110011111111111111001111111111111101;
    wire [5:0] lut_810_select = {
                             in_data[132],
                             in_data[533],
                             in_data[253],
                             in_data[109],
                             in_data[767],
                             in_data[81]};
    
    wire lut_810_out = lut_810_table[lut_810_select];
    
    generate
    if ( USE_REG ) begin : ff_810
        reg   lut_810_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_810_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_810_ff <= lut_810_out;
            end
        end
        
        assign out_data[810] = lut_810_ff;
    end
    else begin : no_ff_810
        assign out_data[810] = lut_810_out;
    end
    endgenerate
    
    
    
    // LUT : 811
    wire [63:0] lut_811_table = 64'b1111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_811_select = {
                             in_data[255],
                             in_data[107],
                             in_data[475],
                             in_data[158],
                             in_data[98],
                             in_data[126]};
    
    wire lut_811_out = lut_811_table[lut_811_select];
    
    generate
    if ( USE_REG ) begin : ff_811
        reg   lut_811_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_811_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_811_ff <= lut_811_out;
            end
        end
        
        assign out_data[811] = lut_811_ff;
    end
    else begin : no_ff_811
        assign out_data[811] = lut_811_out;
    end
    endgenerate
    
    
    
    // LUT : 812
    wire [63:0] lut_812_table = 64'b0000000011010100000011111111111100000000000000001000111110001111;
    wire [5:0] lut_812_select = {
                             in_data[545],
                             in_data[543],
                             in_data[657],
                             in_data[245],
                             in_data[182],
                             in_data[64]};
    
    wire lut_812_out = lut_812_table[lut_812_select];
    
    generate
    if ( USE_REG ) begin : ff_812
        reg   lut_812_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_812_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_812_ff <= lut_812_out;
            end
        end
        
        assign out_data[812] = lut_812_ff;
    end
    else begin : no_ff_812
        assign out_data[812] = lut_812_out;
    end
    endgenerate
    
    
    
    // LUT : 813
    wire [63:0] lut_813_table = 64'b0000010100000000000000000000000001010101000001010101010100000101;
    wire [5:0] lut_813_select = {
                             in_data[650],
                             in_data[254],
                             in_data[247],
                             in_data[556],
                             in_data[252],
                             in_data[175]};
    
    wire lut_813_out = lut_813_table[lut_813_select];
    
    generate
    if ( USE_REG ) begin : ff_813
        reg   lut_813_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_813_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_813_ff <= lut_813_out;
            end
        end
        
        assign out_data[813] = lut_813_ff;
    end
    else begin : no_ff_813
        assign out_data[813] = lut_813_out;
    end
    endgenerate
    
    
    
    // LUT : 814
    wire [63:0] lut_814_table = 64'b0000000000000000001100000011000000000000000000000011000000110000;
    wire [5:0] lut_814_select = {
                             in_data[737],
                             in_data[199],
                             in_data[91],
                             in_data[456],
                             in_data[257],
                             in_data[477]};
    
    wire lut_814_out = lut_814_table[lut_814_select];
    
    generate
    if ( USE_REG ) begin : ff_814
        reg   lut_814_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_814_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_814_ff <= lut_814_out;
            end
        end
        
        assign out_data[814] = lut_814_ff;
    end
    else begin : no_ff_814
        assign out_data[814] = lut_814_out;
    end
    endgenerate
    
    
    
    // LUT : 815
    wire [63:0] lut_815_table = 64'b0000000010000000000000000000000010101010101010101010101010101010;
    wire [5:0] lut_815_select = {
                             in_data[573],
                             in_data[726],
                             in_data[145],
                             in_data[504],
                             in_data[280],
                             in_data[261]};
    
    wire lut_815_out = lut_815_table[lut_815_select];
    
    generate
    if ( USE_REG ) begin : ff_815
        reg   lut_815_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_815_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_815_ff <= lut_815_out;
            end
        end
        
        assign out_data[815] = lut_815_ff;
    end
    else begin : no_ff_815
        assign out_data[815] = lut_815_out;
    end
    endgenerate
    
    
    
    // LUT : 816
    wire [63:0] lut_816_table = 64'b1111111111111111111111111111111011111111111111001111110011001100;
    wire [5:0] lut_816_select = {
                             in_data[212],
                             in_data[68],
                             in_data[523],
                             in_data[11],
                             in_data[304],
                             in_data[647]};
    
    wire lut_816_out = lut_816_table[lut_816_select];
    
    generate
    if ( USE_REG ) begin : ff_816
        reg   lut_816_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_816_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_816_ff <= lut_816_out;
            end
        end
        
        assign out_data[816] = lut_816_ff;
    end
    else begin : no_ff_816
        assign out_data[816] = lut_816_out;
    end
    endgenerate
    
    
    
    // LUT : 817
    wire [63:0] lut_817_table = 64'b1111111100000000010101010000000011111111101010111111111110101010;
    wire [5:0] lut_817_select = {
                             in_data[746],
                             in_data[623],
                             in_data[231],
                             in_data[447],
                             in_data[139],
                             in_data[605]};
    
    wire lut_817_out = lut_817_table[lut_817_select];
    
    generate
    if ( USE_REG ) begin : ff_817
        reg   lut_817_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_817_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_817_ff <= lut_817_out;
            end
        end
        
        assign out_data[817] = lut_817_ff;
    end
    else begin : no_ff_817
        assign out_data[817] = lut_817_out;
    end
    endgenerate
    
    
    
    // LUT : 818
    wire [63:0] lut_818_table = 64'b0000000000000000000011110000111000000000000000000000111100001110;
    wire [5:0] lut_818_select = {
                             in_data[15],
                             in_data[144],
                             in_data[339],
                             in_data[74],
                             in_data[146],
                             in_data[590]};
    
    wire lut_818_out = lut_818_table[lut_818_select];
    
    generate
    if ( USE_REG ) begin : ff_818
        reg   lut_818_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_818_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_818_ff <= lut_818_out;
            end
        end
        
        assign out_data[818] = lut_818_ff;
    end
    else begin : no_ff_818
        assign out_data[818] = lut_818_out;
    end
    endgenerate
    
    
    
    // LUT : 819
    wire [63:0] lut_819_table = 64'b1111111011101110111111101110110011111110111011101111111011101100;
    wire [5:0] lut_819_select = {
                             in_data[752],
                             in_data[292],
                             in_data[312],
                             in_data[423],
                             in_data[400],
                             in_data[404]};
    
    wire lut_819_out = lut_819_table[lut_819_select];
    
    generate
    if ( USE_REG ) begin : ff_819
        reg   lut_819_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_819_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_819_ff <= lut_819_out;
            end
        end
        
        assign out_data[819] = lut_819_ff;
    end
    else begin : no_ff_819
        assign out_data[819] = lut_819_out;
    end
    endgenerate
    
    
    
    // LUT : 820
    wire [63:0] lut_820_table = 64'b0000000000000000000000001010111100000000000000000000000010101011;
    wire [5:0] lut_820_select = {
                             in_data[589],
                             in_data[610],
                             in_data[133],
                             in_data[656],
                             in_data[747],
                             in_data[177]};
    
    wire lut_820_out = lut_820_table[lut_820_select];
    
    generate
    if ( USE_REG ) begin : ff_820
        reg   lut_820_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_820_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_820_ff <= lut_820_out;
            end
        end
        
        assign out_data[820] = lut_820_ff;
    end
    else begin : no_ff_820
        assign out_data[820] = lut_820_out;
    end
    endgenerate
    
    
    
    // LUT : 821
    wire [63:0] lut_821_table = 64'b1111111111111111111110111111111111111011111111111111001111110011;
    wire [5:0] lut_821_select = {
                             in_data[221],
                             in_data[666],
                             in_data[618],
                             in_data[689],
                             in_data[631],
                             in_data[94]};
    
    wire lut_821_out = lut_821_table[lut_821_select];
    
    generate
    if ( USE_REG ) begin : ff_821
        reg   lut_821_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_821_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_821_ff <= lut_821_out;
            end
        end
        
        assign out_data[821] = lut_821_ff;
    end
    else begin : no_ff_821
        assign out_data[821] = lut_821_out;
    end
    endgenerate
    
    
    
    // LUT : 822
    wire [63:0] lut_822_table = 64'b1111111110101010111111110000000010111111101010101111111100000000;
    wire [5:0] lut_822_select = {
                             in_data[51],
                             in_data[662],
                             in_data[348],
                             in_data[364],
                             in_data[205],
                             in_data[653]};
    
    wire lut_822_out = lut_822_table[lut_822_select];
    
    generate
    if ( USE_REG ) begin : ff_822
        reg   lut_822_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_822_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_822_ff <= lut_822_out;
            end
        end
        
        assign out_data[822] = lut_822_ff;
    end
    else begin : no_ff_822
        assign out_data[822] = lut_822_out;
    end
    endgenerate
    
    
    
    // LUT : 823
    wire [63:0] lut_823_table = 64'b1111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_823_select = {
                             in_data[588],
                             in_data[736],
                             in_data[757],
                             in_data[232],
                             in_data[714],
                             in_data[532]};
    
    wire lut_823_out = lut_823_table[lut_823_select];
    
    generate
    if ( USE_REG ) begin : ff_823
        reg   lut_823_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_823_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_823_ff <= lut_823_out;
            end
        end
        
        assign out_data[823] = lut_823_ff;
    end
    else begin : no_ff_823
        assign out_data[823] = lut_823_out;
    end
    endgenerate
    
    
    
    // LUT : 824
    wire [63:0] lut_824_table = 64'b1111111100000111111111110000000011111111000011111111111100000000;
    wire [5:0] lut_824_select = {
                             in_data[774],
                             in_data[687],
                             in_data[289],
                             in_data[164],
                             in_data[478],
                             in_data[89]};
    
    wire lut_824_out = lut_824_table[lut_824_select];
    
    generate
    if ( USE_REG ) begin : ff_824
        reg   lut_824_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_824_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_824_ff <= lut_824_out;
            end
        end
        
        assign out_data[824] = lut_824_ff;
    end
    else begin : no_ff_824
        assign out_data[824] = lut_824_out;
    end
    endgenerate
    
    
    
    // LUT : 825
    wire [63:0] lut_825_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_825_select = {
                             in_data[87],
                             in_data[56],
                             in_data[643],
                             in_data[780],
                             in_data[376],
                             in_data[615]};
    
    wire lut_825_out = lut_825_table[lut_825_select];
    
    generate
    if ( USE_REG ) begin : ff_825
        reg   lut_825_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_825_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_825_ff <= lut_825_out;
            end
        end
        
        assign out_data[825] = lut_825_ff;
    end
    else begin : no_ff_825
        assign out_data[825] = lut_825_out;
    end
    endgenerate
    
    
    
    // LUT : 826
    wire [63:0] lut_826_table = 64'b0101000011111111010100001111111001010000111111110101000011111110;
    wire [5:0] lut_826_select = {
                             in_data[763],
                             in_data[472],
                             in_data[467],
                             in_data[327],
                             in_data[19],
                             in_data[660]};
    
    wire lut_826_out = lut_826_table[lut_826_select];
    
    generate
    if ( USE_REG ) begin : ff_826
        reg   lut_826_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_826_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_826_ff <= lut_826_out;
            end
        end
        
        assign out_data[826] = lut_826_ff;
    end
    else begin : no_ff_826
        assign out_data[826] = lut_826_out;
    end
    endgenerate
    
    
    
    // LUT : 827
    wire [63:0] lut_827_table = 64'b0010101110101011000000111010101100101011101010110000001110101011;
    wire [5:0] lut_827_select = {
                             in_data[783],
                             in_data[512],
                             in_data[272],
                             in_data[235],
                             in_data[554],
                             in_data[101]};
    
    wire lut_827_out = lut_827_table[lut_827_select];
    
    generate
    if ( USE_REG ) begin : ff_827
        reg   lut_827_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_827_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_827_ff <= lut_827_out;
            end
        end
        
        assign out_data[827] = lut_827_ff;
    end
    else begin : no_ff_827
        assign out_data[827] = lut_827_out;
    end
    endgenerate
    
    
    
    // LUT : 828
    wire [63:0] lut_828_table = 64'b0000001010101011000000000010001100000000101110110010000000100011;
    wire [5:0] lut_828_select = {
                             in_data[365],
                             in_data[153],
                             in_data[526],
                             in_data[673],
                             in_data[482],
                             in_data[242]};
    
    wire lut_828_out = lut_828_table[lut_828_select];
    
    generate
    if ( USE_REG ) begin : ff_828
        reg   lut_828_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_828_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_828_ff <= lut_828_out;
            end
        end
        
        assign out_data[828] = lut_828_ff;
    end
    else begin : no_ff_828
        assign out_data[828] = lut_828_out;
    end
    endgenerate
    
    
    
    // LUT : 829
    wire [63:0] lut_829_table = 64'b0011001111111111001100111111111100010001110111010011000111011101;
    wire [5:0] lut_829_select = {
                             in_data[688],
                             in_data[674],
                             in_data[494],
                             in_data[196],
                             in_data[412],
                             in_data[121]};
    
    wire lut_829_out = lut_829_table[lut_829_select];
    
    generate
    if ( USE_REG ) begin : ff_829
        reg   lut_829_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_829_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_829_ff <= lut_829_out;
            end
        end
        
        assign out_data[829] = lut_829_ff;
    end
    else begin : no_ff_829
        assign out_data[829] = lut_829_out;
    end
    endgenerate
    
    
    
    // LUT : 830
    wire [63:0] lut_830_table = 64'b0000001000000010000000100000001000101011001010110010101100101011;
    wire [5:0] lut_830_select = {
                             in_data[637],
                             in_data[39],
                             in_data[755],
                             in_data[381],
                             in_data[149],
                             in_data[385]};
    
    wire lut_830_out = lut_830_table[lut_830_select];
    
    generate
    if ( USE_REG ) begin : ff_830
        reg   lut_830_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_830_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_830_ff <= lut_830_out;
            end
        end
        
        assign out_data[830] = lut_830_ff;
    end
    else begin : no_ff_830
        assign out_data[830] = lut_830_out;
    end
    endgenerate
    
    
    
    // LUT : 831
    wire [63:0] lut_831_table = 64'b0000000000000000000000000000000000001111000011110000111100001111;
    wire [5:0] lut_831_select = {
                             in_data[360],
                             in_data[754],
                             in_data[114],
                             in_data[186],
                             in_data[421],
                             in_data[730]};
    
    wire lut_831_out = lut_831_table[lut_831_select];
    
    generate
    if ( USE_REG ) begin : ff_831
        reg   lut_831_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_831_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_831_ff <= lut_831_out;
            end
        end
        
        assign out_data[831] = lut_831_ff;
    end
    else begin : no_ff_831
        assign out_data[831] = lut_831_out;
    end
    endgenerate
    
    
    
    // LUT : 832
    wire [63:0] lut_832_table = 64'b1101110111011101110111011101110111111111010101011111111101010101;
    wire [5:0] lut_832_select = {
                             in_data[595],
                             in_data[699],
                             in_data[681],
                             in_data[201],
                             in_data[407],
                             in_data[484]};
    
    wire lut_832_out = lut_832_table[lut_832_select];
    
    generate
    if ( USE_REG ) begin : ff_832
        reg   lut_832_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_832_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_832_ff <= lut_832_out;
            end
        end
        
        assign out_data[832] = lut_832_ff;
    end
    else begin : no_ff_832
        assign out_data[832] = lut_832_out;
    end
    endgenerate
    
    
    
    // LUT : 833
    wire [63:0] lut_833_table = 64'b0101000011010100010100001101010101010000110101010101000011010101;
    wire [5:0] lut_833_select = {
                             in_data[78],
                             in_data[120],
                             in_data[440],
                             in_data[632],
                             in_data[246],
                             in_data[540]};
    
    wire lut_833_out = lut_833_table[lut_833_select];
    
    generate
    if ( USE_REG ) begin : ff_833
        reg   lut_833_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_833_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_833_ff <= lut_833_out;
            end
        end
        
        assign out_data[833] = lut_833_ff;
    end
    else begin : no_ff_833
        assign out_data[833] = lut_833_out;
    end
    endgenerate
    
    
    
    // LUT : 834
    wire [63:0] lut_834_table = 64'b1000111100001100100011110000110011101111000011011010111100001101;
    wire [5:0] lut_834_select = {
                             in_data[417],
                             in_data[503],
                             in_data[734],
                             in_data[581],
                             in_data[716],
                             in_data[331]};
    
    wire lut_834_out = lut_834_table[lut_834_select];
    
    generate
    if ( USE_REG ) begin : ff_834
        reg   lut_834_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_834_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_834_ff <= lut_834_out;
            end
        end
        
        assign out_data[834] = lut_834_ff;
    end
    else begin : no_ff_834
        assign out_data[834] = lut_834_out;
    end
    endgenerate
    
    
    
    // LUT : 835
    wire [63:0] lut_835_table = 64'b0101010100000011010100010000001101010001000000110101000100000011;
    wire [5:0] lut_835_select = {
                             in_data[137],
                             in_data[36],
                             in_data[654],
                             in_data[382],
                             in_data[413],
                             in_data[619]};
    
    wire lut_835_out = lut_835_table[lut_835_select];
    
    generate
    if ( USE_REG ) begin : ff_835
        reg   lut_835_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_835_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_835_ff <= lut_835_out;
            end
        end
        
        assign out_data[835] = lut_835_ff;
    end
    else begin : no_ff_835
        assign out_data[835] = lut_835_out;
    end
    endgenerate
    
    
    
    // LUT : 836
    wire [63:0] lut_836_table = 64'b0011000011111111011000001111111100000000111100001100000011111100;
    wire [5:0] lut_836_select = {
                             in_data[191],
                             in_data[713],
                             in_data[667],
                             in_data[192],
                             in_data[359],
                             in_data[63]};
    
    wire lut_836_out = lut_836_table[lut_836_select];
    
    generate
    if ( USE_REG ) begin : ff_836
        reg   lut_836_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_836_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_836_ff <= lut_836_out;
            end
        end
        
        assign out_data[836] = lut_836_ff;
    end
    else begin : no_ff_836
        assign out_data[836] = lut_836_out;
    end
    endgenerate
    
    
    
    // LUT : 837
    wire [63:0] lut_837_table = 64'b0011111100111011001111110011101100110011001100110011001100110011;
    wire [5:0] lut_837_select = {
                             in_data[181],
                             in_data[765],
                             in_data[305],
                             in_data[372],
                             in_data[492],
                             in_data[227]};
    
    wire lut_837_out = lut_837_table[lut_837_select];
    
    generate
    if ( USE_REG ) begin : ff_837
        reg   lut_837_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_837_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_837_ff <= lut_837_out;
            end
        end
        
        assign out_data[837] = lut_837_ff;
    end
    else begin : no_ff_837
        assign out_data[837] = lut_837_out;
    end
    endgenerate
    
    
    
    // LUT : 838
    wire [63:0] lut_838_table = 64'b0000000001010101000001001101111100000000010101010000010011011111;
    wire [5:0] lut_838_select = {
                             in_data[9],
                             in_data[441],
                             in_data[263],
                             in_data[310],
                             in_data[202],
                             in_data[715]};
    
    wire lut_838_out = lut_838_table[lut_838_select];
    
    generate
    if ( USE_REG ) begin : ff_838
        reg   lut_838_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_838_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_838_ff <= lut_838_out;
            end
        end
        
        assign out_data[838] = lut_838_ff;
    end
    else begin : no_ff_838
        assign out_data[838] = lut_838_out;
    end
    endgenerate
    
    
    
    // LUT : 839
    wire [63:0] lut_839_table = 64'b0101010001010000010101000101000001010100010101010101010001010101;
    wire [5:0] lut_839_select = {
                             in_data[313],
                             in_data[62],
                             in_data[663],
                             in_data[629],
                             in_data[45],
                             in_data[301]};
    
    wire lut_839_out = lut_839_table[lut_839_select];
    
    generate
    if ( USE_REG ) begin : ff_839
        reg   lut_839_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_839_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_839_ff <= lut_839_out;
            end
        end
        
        assign out_data[839] = lut_839_ff;
    end
    else begin : no_ff_839
        assign out_data[839] = lut_839_out;
    end
    endgenerate
    
    
    
    // LUT : 840
    wire [63:0] lut_840_table = 64'b0101010101010101000000000000000000000101000001010000010000000000;
    wire [5:0] lut_840_select = {
                             in_data[179],
                             in_data[491],
                             in_data[106],
                             in_data[593],
                             in_data[115],
                             in_data[277]};
    
    wire lut_840_out = lut_840_table[lut_840_select];
    
    generate
    if ( USE_REG ) begin : ff_840
        reg   lut_840_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_840_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_840_ff <= lut_840_out;
            end
        end
        
        assign out_data[840] = lut_840_ff;
    end
    else begin : no_ff_840
        assign out_data[840] = lut_840_out;
    end
    endgenerate
    
    
    
    // LUT : 841
    wire [63:0] lut_841_table = 64'b0100010101010101000001010001110101000101010001010000010100000101;
    wire [5:0] lut_841_select = {
                             in_data[185],
                             in_data[4],
                             in_data[251],
                             in_data[134],
                             in_data[275],
                             in_data[411]};
    
    wire lut_841_out = lut_841_table[lut_841_select];
    
    generate
    if ( USE_REG ) begin : ff_841
        reg   lut_841_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_841_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_841_ff <= lut_841_out;
            end
        end
        
        assign out_data[841] = lut_841_ff;
    end
    else begin : no_ff_841
        assign out_data[841] = lut_841_out;
    end
    endgenerate
    
    
    
    // LUT : 842
    wire [63:0] lut_842_table = 64'b0000000000000000111111111111111100000000000000001000000011000100;
    wire [5:0] lut_842_select = {
                             in_data[522],
                             in_data[594],
                             in_data[587],
                             in_data[93],
                             in_data[165],
                             in_data[7]};
    
    wire lut_842_out = lut_842_table[lut_842_select];
    
    generate
    if ( USE_REG ) begin : ff_842
        reg   lut_842_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_842_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_842_ff <= lut_842_out;
            end
        end
        
        assign out_data[842] = lut_842_ff;
    end
    else begin : no_ff_842
        assign out_data[842] = lut_842_out;
    end
    endgenerate
    
    
    
    // LUT : 843
    wire [63:0] lut_843_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_843_select = {
                             in_data[358],
                             in_data[583],
                             in_data[749],
                             in_data[596],
                             in_data[97],
                             in_data[18]};
    
    wire lut_843_out = lut_843_table[lut_843_select];
    
    generate
    if ( USE_REG ) begin : ff_843
        reg   lut_843_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_843_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_843_ff <= lut_843_out;
            end
        end
        
        assign out_data[843] = lut_843_ff;
    end
    else begin : no_ff_843
        assign out_data[843] = lut_843_out;
    end
    endgenerate
    
    
    
    // LUT : 844
    wire [63:0] lut_844_table = 64'b0011001100110011001100110011001100000011000000110000111100001111;
    wire [5:0] lut_844_select = {
                             in_data[680],
                             in_data[129],
                             in_data[693],
                             in_data[462],
                             in_data[189],
                             in_data[727]};
    
    wire lut_844_out = lut_844_table[lut_844_select];
    
    generate
    if ( USE_REG ) begin : ff_844
        reg   lut_844_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_844_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_844_ff <= lut_844_out;
            end
        end
        
        assign out_data[844] = lut_844_ff;
    end
    else begin : no_ff_844
        assign out_data[844] = lut_844_out;
    end
    endgenerate
    
    
    
    // LUT : 845
    wire [63:0] lut_845_table = 64'b1100111111001111110011111100111111001111110011111100111111001111;
    wire [5:0] lut_845_select = {
                             in_data[26],
                             in_data[334],
                             in_data[25],
                             in_data[464],
                             in_data[745],
                             in_data[342]};
    
    wire lut_845_out = lut_845_table[lut_845_select];
    
    generate
    if ( USE_REG ) begin : ff_845
        reg   lut_845_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_845_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_845_ff <= lut_845_out;
            end
        end
        
        assign out_data[845] = lut_845_ff;
    end
    else begin : no_ff_845
        assign out_data[845] = lut_845_out;
    end
    endgenerate
    
    
    
    // LUT : 846
    wire [63:0] lut_846_table = 64'b0000000000000000001000101111111100000000000000000000001111111111;
    wire [5:0] lut_846_select = {
                             in_data[766],
                             in_data[518],
                             in_data[238],
                             in_data[57],
                             in_data[640],
                             in_data[560]};
    
    wire lut_846_out = lut_846_table[lut_846_select];
    
    generate
    if ( USE_REG ) begin : ff_846
        reg   lut_846_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_846_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_846_ff <= lut_846_out;
            end
        end
        
        assign out_data[846] = lut_846_ff;
    end
    else begin : no_ff_846
        assign out_data[846] = lut_846_out;
    end
    endgenerate
    
    
    
    // LUT : 847
    wire [63:0] lut_847_table = 64'b0000000011110000111100001111111001000000111100001100000011111100;
    wire [5:0] lut_847_select = {
                             in_data[652],
                             in_data[524],
                             in_data[102],
                             in_data[268],
                             in_data[592],
                             in_data[113]};
    
    wire lut_847_out = lut_847_table[lut_847_select];
    
    generate
    if ( USE_REG ) begin : ff_847
        reg   lut_847_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_847_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_847_ff <= lut_847_out;
            end
        end
        
        assign out_data[847] = lut_847_ff;
    end
    else begin : no_ff_847
        assign out_data[847] = lut_847_out;
    end
    endgenerate
    
    
    
    // LUT : 848
    wire [63:0] lut_848_table = 64'b0000000000000000000000000000000000000000000000000000000001010101;
    wire [5:0] lut_848_select = {
                             in_data[222],
                             in_data[682],
                             in_data[206],
                             in_data[728],
                             in_data[772],
                             in_data[579]};
    
    wire lut_848_out = lut_848_table[lut_848_select];
    
    generate
    if ( USE_REG ) begin : ff_848
        reg   lut_848_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_848_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_848_ff <= lut_848_out;
            end
        end
        
        assign out_data[848] = lut_848_ff;
    end
    else begin : no_ff_848
        assign out_data[848] = lut_848_out;
    end
    endgenerate
    
    
    
    // LUT : 849
    wire [63:0] lut_849_table = 64'b0000111100001111000010100000101100001111000011110000101100001010;
    wire [5:0] lut_849_select = {
                             in_data[698],
                             in_data[549],
                             in_data[77],
                             in_data[386],
                             in_data[770],
                             in_data[602]};
    
    wire lut_849_out = lut_849_table[lut_849_select];
    
    generate
    if ( USE_REG ) begin : ff_849
        reg   lut_849_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_849_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_849_ff <= lut_849_out;
            end
        end
        
        assign out_data[849] = lut_849_ff;
    end
    else begin : no_ff_849
        assign out_data[849] = lut_849_out;
    end
    endgenerate
    
    
    
    // LUT : 850
    wire [63:0] lut_850_table = 64'b0101010101010101010101010101010101010101010101010101010101010101;
    wire [5:0] lut_850_select = {
                             in_data[154],
                             in_data[168],
                             in_data[762],
                             in_data[642],
                             in_data[328],
                             in_data[598]};
    
    wire lut_850_out = lut_850_table[lut_850_select];
    
    generate
    if ( USE_REG ) begin : ff_850
        reg   lut_850_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_850_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_850_ff <= lut_850_out;
            end
        end
        
        assign out_data[850] = lut_850_ff;
    end
    else begin : no_ff_850
        assign out_data[850] = lut_850_out;
    end
    endgenerate
    
    
    
    // LUT : 851
    wire [63:0] lut_851_table = 64'b1111111111111111000011000000110011111111111111110000110000001100;
    wire [5:0] lut_851_select = {
                             in_data[340],
                             in_data[599],
                             in_data[49],
                             in_data[686],
                             in_data[442],
                             in_data[646]};
    
    wire lut_851_out = lut_851_table[lut_851_select];
    
    generate
    if ( USE_REG ) begin : ff_851
        reg   lut_851_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_851_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_851_ff <= lut_851_out;
            end
        end
        
        assign out_data[851] = lut_851_ff;
    end
    else begin : no_ff_851
        assign out_data[851] = lut_851_out;
    end
    endgenerate
    
    
    
    // LUT : 852
    wire [63:0] lut_852_table = 64'b1110111100001111111011111010111111001100000011001010111110001111;
    wire [5:0] lut_852_select = {
                             in_data[66],
                             in_data[216],
                             in_data[537],
                             in_data[264],
                             in_data[466],
                             in_data[634]};
    
    wire lut_852_out = lut_852_table[lut_852_select];
    
    generate
    if ( USE_REG ) begin : ff_852
        reg   lut_852_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_852_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_852_ff <= lut_852_out;
            end
        end
        
        assign out_data[852] = lut_852_ff;
    end
    else begin : no_ff_852
        assign out_data[852] = lut_852_out;
    end
    endgenerate
    
    
    
    // LUT : 853
    wire [63:0] lut_853_table = 64'b1111111111111111111011101110111011101110111011101110101011101010;
    wire [5:0] lut_853_select = {
                             in_data[237],
                             in_data[748],
                             in_data[42],
                             in_data[1],
                             in_data[433],
                             in_data[487]};
    
    wire lut_853_out = lut_853_table[lut_853_select];
    
    generate
    if ( USE_REG ) begin : ff_853
        reg   lut_853_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_853_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_853_ff <= lut_853_out;
            end
        end
        
        assign out_data[853] = lut_853_ff;
    end
    else begin : no_ff_853
        assign out_data[853] = lut_853_out;
    end
    endgenerate
    
    
    
    // LUT : 854
    wire [63:0] lut_854_table = 64'b1100110011001100111011101110111011101110111011101111111111101111;
    wire [5:0] lut_854_select = {
                             in_data[178],
                             in_data[155],
                             in_data[40],
                             in_data[641],
                             in_data[103],
                             in_data[694]};
    
    wire lut_854_out = lut_854_table[lut_854_select];
    
    generate
    if ( USE_REG ) begin : ff_854
        reg   lut_854_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_854_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_854_ff <= lut_854_out;
            end
        end
        
        assign out_data[854] = lut_854_ff;
    end
    else begin : no_ff_854
        assign out_data[854] = lut_854_out;
    end
    endgenerate
    
    
    
    // LUT : 855
    wire [63:0] lut_855_table = 64'b1010111001010000101011110101000010101110010100001010111101010000;
    wire [5:0] lut_855_select = {
                             in_data[281],
                             in_data[706],
                             in_data[569],
                             in_data[431],
                             in_data[124],
                             in_data[567]};
    
    wire lut_855_out = lut_855_table[lut_855_select];
    
    generate
    if ( USE_REG ) begin : ff_855
        reg   lut_855_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_855_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_855_ff <= lut_855_out;
            end
        end
        
        assign out_data[855] = lut_855_ff;
    end
    else begin : no_ff_855
        assign out_data[855] = lut_855_out;
    end
    endgenerate
    
    
    
    // LUT : 856
    wire [63:0] lut_856_table = 64'b1010101010101010101010101010101011111101111110101111110111101010;
    wire [5:0] lut_856_select = {
                             in_data[461],
                             in_data[675],
                             in_data[127],
                             in_data[719],
                             in_data[709],
                             in_data[353]};
    
    wire lut_856_out = lut_856_table[lut_856_select];
    
    generate
    if ( USE_REG ) begin : ff_856
        reg   lut_856_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_856_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_856_ff <= lut_856_out;
            end
        end
        
        assign out_data[856] = lut_856_ff;
    end
    else begin : no_ff_856
        assign out_data[856] = lut_856_out;
    end
    endgenerate
    
    
    
    // LUT : 857
    wire [63:0] lut_857_table = 64'b1111111100000000111111110000000011111111111111111111111111111111;
    wire [5:0] lut_857_select = {
                             in_data[459],
                             in_data[711],
                             in_data[256],
                             in_data[616],
                             in_data[17],
                             in_data[197]};
    
    wire lut_857_out = lut_857_table[lut_857_select];
    
    generate
    if ( USE_REG ) begin : ff_857
        reg   lut_857_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_857_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_857_ff <= lut_857_out;
            end
        end
        
        assign out_data[857] = lut_857_ff;
    end
    else begin : no_ff_857
        assign out_data[857] = lut_857_out;
    end
    endgenerate
    
    
    
    // LUT : 858
    wire [63:0] lut_858_table = 64'b1110111111001111110011111100111111001110110011101100111111001110;
    wire [5:0] lut_858_select = {
                             in_data[528],
                             in_data[722],
                             in_data[513],
                             in_data[183],
                             in_data[233],
                             in_data[240]};
    
    wire lut_858_out = lut_858_table[lut_858_select];
    
    generate
    if ( USE_REG ) begin : ff_858
        reg   lut_858_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_858_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_858_ff <= lut_858_out;
            end
        end
        
        assign out_data[858] = lut_858_ff;
    end
    else begin : no_ff_858
        assign out_data[858] = lut_858_out;
    end
    endgenerate
    
    
    
    // LUT : 859
    wire [63:0] lut_859_table = 64'b1010000010000000111111111111101010101010101000001111111111111010;
    wire [5:0] lut_859_select = {
                             in_data[279],
                             in_data[314],
                             in_data[95],
                             in_data[539],
                             in_data[138],
                             in_data[152]};
    
    wire lut_859_out = lut_859_table[lut_859_select];
    
    generate
    if ( USE_REG ) begin : ff_859
        reg   lut_859_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_859_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_859_ff <= lut_859_out;
            end
        end
        
        assign out_data[859] = lut_859_ff;
    end
    else begin : no_ff_859
        assign out_data[859] = lut_859_out;
    end
    endgenerate
    
    
    
    // LUT : 860
    wire [63:0] lut_860_table = 64'b0010001000100010001000100010001010111011101110111011101110111011;
    wire [5:0] lut_860_select = {
                             in_data[718],
                             in_data[782],
                             in_data[561],
                             in_data[739],
                             in_data[457],
                             in_data[525]};
    
    wire lut_860_out = lut_860_table[lut_860_select];
    
    generate
    if ( USE_REG ) begin : ff_860
        reg   lut_860_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_860_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_860_ff <= lut_860_out;
            end
        end
        
        assign out_data[860] = lut_860_ff;
    end
    else begin : no_ff_860
        assign out_data[860] = lut_860_out;
    end
    endgenerate
    
    
    
    // LUT : 861
    wire [63:0] lut_861_table = 64'b0100010000000000010100000011000001010100001001000101010101110111;
    wire [5:0] lut_861_select = {
                             in_data[721],
                             in_data[329],
                             in_data[401],
                             in_data[147],
                             in_data[355],
                             in_data[468]};
    
    wire lut_861_out = lut_861_table[lut_861_select];
    
    generate
    if ( USE_REG ) begin : ff_861
        reg   lut_861_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_861_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_861_ff <= lut_861_out;
            end
        end
        
        assign out_data[861] = lut_861_ff;
    end
    else begin : no_ff_861
        assign out_data[861] = lut_861_out;
    end
    endgenerate
    
    
    
    // LUT : 862
    wire [63:0] lut_862_table = 64'b1111111100101100111111110000110011111111001011001111111100100100;
    wire [5:0] lut_862_select = {
                             in_data[308],
                             in_data[529],
                             in_data[288],
                             in_data[550],
                             in_data[295],
                             in_data[430]};
    
    wire lut_862_out = lut_862_table[lut_862_select];
    
    generate
    if ( USE_REG ) begin : ff_862
        reg   lut_862_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_862_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_862_ff <= lut_862_out;
            end
        end
        
        assign out_data[862] = lut_862_ff;
    end
    else begin : no_ff_862
        assign out_data[862] = lut_862_out;
    end
    endgenerate
    
    
    
    // LUT : 863
    wire [63:0] lut_863_table = 64'b1101111111111111010101010101010101010101111111110000010101010101;
    wire [5:0] lut_863_select = {
                             in_data[282],
                             in_data[105],
                             in_data[248],
                             in_data[363],
                             in_data[37],
                             in_data[542]};
    
    wire lut_863_out = lut_863_table[lut_863_select];
    
    generate
    if ( USE_REG ) begin : ff_863
        reg   lut_863_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_863_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_863_ff <= lut_863_out;
            end
        end
        
        assign out_data[863] = lut_863_ff;
    end
    else begin : no_ff_863
        assign out_data[863] = lut_863_out;
    end
    endgenerate
    
    
    
    // LUT : 864
    wire [63:0] lut_864_table = 64'b1010000010100000111101010101010100000000000000000001010100000101;
    wire [5:0] lut_864_select = {
                             in_data[445],
                             in_data[69],
                             in_data[530],
                             in_data[501],
                             in_data[725],
                             in_data[572]};
    
    wire lut_864_out = lut_864_table[lut_864_select];
    
    generate
    if ( USE_REG ) begin : ff_864
        reg   lut_864_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_864_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_864_ff <= lut_864_out;
            end
        end
        
        assign out_data[864] = lut_864_ff;
    end
    else begin : no_ff_864
        assign out_data[864] = lut_864_out;
    end
    endgenerate
    
    
    
    // LUT : 865
    wire [63:0] lut_865_table = 64'b0011001100110011001100110011001100000000000000110000000000000011;
    wire [5:0] lut_865_select = {
                             in_data[565],
                             in_data[35],
                             in_data[750],
                             in_data[744],
                             in_data[303],
                             in_data[775]};
    
    wire lut_865_out = lut_865_table[lut_865_select];
    
    generate
    if ( USE_REG ) begin : ff_865
        reg   lut_865_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_865_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_865_ff <= lut_865_out;
            end
        end
        
        assign out_data[865] = lut_865_ff;
    end
    else begin : no_ff_865
        assign out_data[865] = lut_865_out;
    end
    endgenerate
    
    
    
    // LUT : 866
    wire [63:0] lut_866_table = 64'b1010101010101010101010101010111010101010101010101010101010101010;
    wire [5:0] lut_866_select = {
                             in_data[214],
                             in_data[639],
                             in_data[270],
                             in_data[695],
                             in_data[638],
                             in_data[626]};
    
    wire lut_866_out = lut_866_table[lut_866_select];
    
    generate
    if ( USE_REG ) begin : ff_866
        reg   lut_866_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_866_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_866_ff <= lut_866_out;
            end
        end
        
        assign out_data[866] = lut_866_ff;
    end
    else begin : no_ff_866
        assign out_data[866] = lut_866_out;
    end
    endgenerate
    
    
    
    // LUT : 867
    wire [63:0] lut_867_table = 64'b1111111111111111111110001111100011111111111111111111100011100000;
    wire [5:0] lut_867_select = {
                             in_data[769],
                             in_data[160],
                             in_data[760],
                             in_data[521],
                             in_data[204],
                             in_data[187]};
    
    wire lut_867_out = lut_867_table[lut_867_select];
    
    generate
    if ( USE_REG ) begin : ff_867
        reg   lut_867_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_867_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_867_ff <= lut_867_out;
            end
        end
        
        assign out_data[867] = lut_867_ff;
    end
    else begin : no_ff_867
        assign out_data[867] = lut_867_out;
    end
    endgenerate
    
    
    
    // LUT : 868
    wire [63:0] lut_868_table = 64'b0111011100000001111111110000000001010101010101000101010101010101;
    wire [5:0] lut_868_select = {
                             in_data[243],
                             in_data[29],
                             in_data[357],
                             in_data[298],
                             in_data[516],
                             in_data[347]};
    
    wire lut_868_out = lut_868_table[lut_868_select];
    
    generate
    if ( USE_REG ) begin : ff_868
        reg   lut_868_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_868_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_868_ff <= lut_868_out;
            end
        end
        
        assign out_data[868] = lut_868_ff;
    end
    else begin : no_ff_868
        assign out_data[868] = lut_868_out;
    end
    endgenerate
    
    
    
    // LUT : 869
    wire [63:0] lut_869_table = 64'b1111111111111111111111111111111111110000111000001111000011010000;
    wire [5:0] lut_869_select = {
                             in_data[297],
                             in_data[283],
                             in_data[117],
                             in_data[259],
                             in_data[741],
                             in_data[23]};
    
    wire lut_869_out = lut_869_table[lut_869_select];
    
    generate
    if ( USE_REG ) begin : ff_869
        reg   lut_869_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_869_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_869_ff <= lut_869_out;
            end
        end
        
        assign out_data[869] = lut_869_ff;
    end
    else begin : no_ff_869
        assign out_data[869] = lut_869_out;
    end
    endgenerate
    
    
    
    // LUT : 870
    wire [63:0] lut_870_table = 64'b0000111100101111000011100000101001010101010101010001000000000000;
    wire [5:0] lut_870_select = {
                             in_data[493],
                             in_data[296],
                             in_data[648],
                             in_data[96],
                             in_data[148],
                             in_data[354]};
    
    wire lut_870_out = lut_870_table[lut_870_select];
    
    generate
    if ( USE_REG ) begin : ff_870
        reg   lut_870_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_870_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_870_ff <= lut_870_out;
            end
        end
        
        assign out_data[870] = lut_870_ff;
    end
    else begin : no_ff_870
        assign out_data[870] = lut_870_out;
    end
    endgenerate
    
    
    
    // LUT : 871
    wire [63:0] lut_871_table = 64'b1111111111111111111111111101111111111111111111111100110011001100;
    wire [5:0] lut_871_select = {
                             in_data[510],
                             in_data[267],
                             in_data[474],
                             in_data[20],
                             in_data[564],
                             in_data[452]};
    
    wire lut_871_out = lut_871_table[lut_871_select];
    
    generate
    if ( USE_REG ) begin : ff_871
        reg   lut_871_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_871_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_871_ff <= lut_871_out;
            end
        end
        
        assign out_data[871] = lut_871_ff;
    end
    else begin : no_ff_871
        assign out_data[871] = lut_871_out;
    end
    endgenerate
    
    
    
    // LUT : 872
    wire [63:0] lut_872_table = 64'b1111111111111111111111111111111111111111111111110000000011110000;
    wire [5:0] lut_872_select = {
                             in_data[351],
                             in_data[325],
                             in_data[90],
                             in_data[370],
                             in_data[28],
                             in_data[751]};
    
    wire lut_872_out = lut_872_table[lut_872_select];
    
    generate
    if ( USE_REG ) begin : ff_872
        reg   lut_872_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_872_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_872_ff <= lut_872_out;
            end
        end
        
        assign out_data[872] = lut_872_ff;
    end
    else begin : no_ff_872
        assign out_data[872] = lut_872_out;
    end
    endgenerate
    
    
    
    // LUT : 873
    wire [63:0] lut_873_table = 64'b0011001100110011000100010001000000110011001100110011001100110011;
    wire [5:0] lut_873_select = {
                             in_data[388],
                             in_data[435],
                             in_data[125],
                             in_data[630],
                             in_data[317],
                             in_data[661]};
    
    wire lut_873_out = lut_873_table[lut_873_select];
    
    generate
    if ( USE_REG ) begin : ff_873
        reg   lut_873_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_873_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_873_ff <= lut_873_out;
            end
        end
        
        assign out_data[873] = lut_873_ff;
    end
    else begin : no_ff_873
        assign out_data[873] = lut_873_out;
    end
    endgenerate
    
    
    
    // LUT : 874
    wire [63:0] lut_874_table = 64'b0000110000000000001011111111111111000000111100001011111111111111;
    wire [5:0] lut_874_select = {
                             in_data[489],
                             in_data[207],
                             in_data[321],
                             in_data[568],
                             in_data[415],
                             in_data[781]};
    
    wire lut_874_out = lut_874_table[lut_874_select];
    
    generate
    if ( USE_REG ) begin : ff_874
        reg   lut_874_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_874_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_874_ff <= lut_874_out;
            end
        end
        
        assign out_data[874] = lut_874_ff;
    end
    else begin : no_ff_874
        assign out_data[874] = lut_874_out;
    end
    endgenerate
    
    
    
    // LUT : 875
    wire [63:0] lut_875_table = 64'b0100000001010000111111001111111011010000110100001111110011111110;
    wire [5:0] lut_875_select = {
                             in_data[384],
                             in_data[239],
                             in_data[773],
                             in_data[511],
                             in_data[375],
                             in_data[379]};
    
    wire lut_875_out = lut_875_table[lut_875_select];
    
    generate
    if ( USE_REG ) begin : ff_875
        reg   lut_875_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_875_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_875_ff <= lut_875_out;
            end
        end
        
        assign out_data[875] = lut_875_ff;
    end
    else begin : no_ff_875
        assign out_data[875] = lut_875_out;
    end
    endgenerate
    
    
    
    // LUT : 876
    wire [63:0] lut_876_table = 64'b1111111110111010111111111010101011111111101111111111111110111010;
    wire [5:0] lut_876_select = {
                             in_data[43],
                             in_data[586],
                             in_data[424],
                             in_data[209],
                             in_data[32],
                             in_data[104]};
    
    wire lut_876_out = lut_876_table[lut_876_select];
    
    generate
    if ( USE_REG ) begin : ff_876
        reg   lut_876_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_876_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_876_ff <= lut_876_out;
            end
        end
        
        assign out_data[876] = lut_876_ff;
    end
    else begin : no_ff_876
        assign out_data[876] = lut_876_out;
    end
    endgenerate
    
    
    
    // LUT : 877
    wire [63:0] lut_877_table = 64'b1010101011111111101010101111111110101010111111111010101011111111;
    wire [5:0] lut_877_select = {
                             in_data[169],
                             in_data[731],
                             in_data[203],
                             in_data[41],
                             in_data[21],
                             in_data[585]};
    
    wire lut_877_out = lut_877_table[lut_877_select];
    
    generate
    if ( USE_REG ) begin : ff_877
        reg   lut_877_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_877_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_877_ff <= lut_877_out;
            end
        end
        
        assign out_data[877] = lut_877_ff;
    end
    else begin : no_ff_877
        assign out_data[877] = lut_877_out;
    end
    endgenerate
    
    
    
    // LUT : 878
    wire [63:0] lut_878_table = 64'b0100010001000100110111011100110001000100010001001101110011001100;
    wire [5:0] lut_878_select = {
                             in_data[198],
                             in_data[458],
                             in_data[38],
                             in_data[278],
                             in_data[436],
                             in_data[692]};
    
    wire lut_878_out = lut_878_table[lut_878_select];
    
    generate
    if ( USE_REG ) begin : ff_878
        reg   lut_878_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_878_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_878_ff <= lut_878_out;
            end
        end
        
        assign out_data[878] = lut_878_ff;
    end
    else begin : no_ff_878
        assign out_data[878] = lut_878_out;
    end
    endgenerate
    
    
    
    // LUT : 879
    wire [63:0] lut_879_table = 64'b0011001100110011101100111011001100110011001100110010001100110011;
    wire [5:0] lut_879_select = {
                             in_data[368],
                             in_data[284],
                             in_data[505],
                             in_data[470],
                             in_data[553],
                             in_data[776]};
    
    wire lut_879_out = lut_879_table[lut_879_select];
    
    generate
    if ( USE_REG ) begin : ff_879
        reg   lut_879_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_879_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_879_ff <= lut_879_out;
            end
        end
        
        assign out_data[879] = lut_879_ff;
    end
    else begin : no_ff_879
        assign out_data[879] = lut_879_out;
    end
    endgenerate
    
    
    
    // LUT : 880
    wire [63:0] lut_880_table = 64'b1111111101001010111111110101111111011010000010101111111101011010;
    wire [5:0] lut_880_select = {
                             in_data[70],
                             in_data[606],
                             in_data[249],
                             in_data[241],
                             in_data[343],
                             in_data[157]};
    
    wire lut_880_out = lut_880_table[lut_880_select];
    
    generate
    if ( USE_REG ) begin : ff_880
        reg   lut_880_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_880_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_880_ff <= lut_880_out;
            end
        end
        
        assign out_data[880] = lut_880_ff;
    end
    else begin : no_ff_880
        assign out_data[880] = lut_880_out;
    end
    endgenerate
    
    
    
    // LUT : 881
    wire [63:0] lut_881_table = 64'b1111111111101110111111111110111001110101000001000111000000000000;
    wire [5:0] lut_881_select = {
                             in_data[519],
                             in_data[777],
                             in_data[396],
                             in_data[409],
                             in_data[580],
                             in_data[374]};
    
    wire lut_881_out = lut_881_table[lut_881_select];
    
    generate
    if ( USE_REG ) begin : ff_881
        reg   lut_881_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_881_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_881_ff <= lut_881_out;
            end
        end
        
        assign out_data[881] = lut_881_ff;
    end
    else begin : no_ff_881
        assign out_data[881] = lut_881_out;
    end
    endgenerate
    
    
    
    // LUT : 882
    wire [63:0] lut_882_table = 64'b1100110011001100110011001100110011111111111111111111111111111110;
    wire [5:0] lut_882_select = {
                             in_data[742],
                             in_data[108],
                             in_data[422],
                             in_data[6],
                             in_data[99],
                             in_data[72]};
    
    wire lut_882_out = lut_882_table[lut_882_select];
    
    generate
    if ( USE_REG ) begin : ff_882
        reg   lut_882_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_882_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_882_ff <= lut_882_out;
            end
        end
        
        assign out_data[882] = lut_882_ff;
    end
    else begin : no_ff_882
        assign out_data[882] = lut_882_out;
    end
    endgenerate
    
    
    
    // LUT : 883
    wire [63:0] lut_883_table = 64'b0000110000001100000011000000110000001000000011000000110000001100;
    wire [5:0] lut_883_select = {
                             in_data[80],
                             in_data[258],
                             in_data[119],
                             in_data[527],
                             in_data[383],
                             in_data[450]};
    
    wire lut_883_out = lut_883_table[lut_883_select];
    
    generate
    if ( USE_REG ) begin : ff_883
        reg   lut_883_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_883_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_883_ff <= lut_883_out;
            end
        end
        
        assign out_data[883] = lut_883_ff;
    end
    else begin : no_ff_883
        assign out_data[883] = lut_883_out;
    end
    endgenerate
    
    
    
    // LUT : 884
    wire [63:0] lut_884_table = 64'b1111111111110111111100101111000011101110000000101110000001110000;
    wire [5:0] lut_884_select = {
                             in_data[577],
                             in_data[576],
                             in_data[575],
                             in_data[548],
                             in_data[271],
                             in_data[600]};
    
    wire lut_884_out = lut_884_table[lut_884_select];
    
    generate
    if ( USE_REG ) begin : ff_884
        reg   lut_884_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_884_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_884_ff <= lut_884_out;
            end
        end
        
        assign out_data[884] = lut_884_ff;
    end
    else begin : no_ff_884
        assign out_data[884] = lut_884_out;
    end
    endgenerate
    
    
    
    // LUT : 885
    wire [63:0] lut_885_table = 64'b1111111111111110111111001111110011111111111111111111010011110000;
    wire [5:0] lut_885_select = {
                             in_data[659],
                             in_data[176],
                             in_data[48],
                             in_data[514],
                             in_data[517],
                             in_data[167]};
    
    wire lut_885_out = lut_885_table[lut_885_select];
    
    generate
    if ( USE_REG ) begin : ff_885
        reg   lut_885_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_885_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_885_ff <= lut_885_out;
            end
        end
        
        assign out_data[885] = lut_885_ff;
    end
    else begin : no_ff_885
        assign out_data[885] = lut_885_out;
    end
    endgenerate
    
    
    
    // LUT : 886
    wire [63:0] lut_886_table = 64'b1111111111001100111111001100110011111111111111111111110011111100;
    wire [5:0] lut_886_select = {
                             in_data[162],
                             in_data[555],
                             in_data[679],
                             in_data[582],
                             in_data[500],
                             in_data[0]};
    
    wire lut_886_out = lut_886_table[lut_886_select];
    
    generate
    if ( USE_REG ) begin : ff_886
        reg   lut_886_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_886_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_886_ff <= lut_886_out;
            end
        end
        
        assign out_data[886] = lut_886_ff;
    end
    else begin : no_ff_886
        assign out_data[886] = lut_886_out;
    end
    endgenerate
    
    
    
    // LUT : 887
    wire [63:0] lut_887_table = 64'b0001010100010101000100010000000101010101000100010001000100010001;
    wire [5:0] lut_887_select = {
                             in_data[55],
                             in_data[768],
                             in_data[559],
                             in_data[142],
                             in_data[488],
                             in_data[79]};
    
    wire lut_887_out = lut_887_table[lut_887_select];
    
    generate
    if ( USE_REG ) begin : ff_887
        reg   lut_887_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_887_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_887_ff <= lut_887_out;
            end
        end
        
        assign out_data[887] = lut_887_ff;
    end
    else begin : no_ff_887
        assign out_data[887] = lut_887_out;
    end
    endgenerate
    
    
    
    // LUT : 888
    wire [63:0] lut_888_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_888_select = {
                             in_data[378],
                             in_data[31],
                             in_data[344],
                             in_data[46],
                             in_data[10],
                             in_data[307]};
    
    wire lut_888_out = lut_888_table[lut_888_select];
    
    generate
    if ( USE_REG ) begin : ff_888
        reg   lut_888_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_888_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_888_ff <= lut_888_out;
            end
        end
        
        assign out_data[888] = lut_888_ff;
    end
    else begin : no_ff_888
        assign out_data[888] = lut_888_out;
    end
    endgenerate
    
    
    
    // LUT : 889
    wire [63:0] lut_889_table = 64'b0010001000100010001000100010001000100010001000100010001000100010;
    wire [5:0] lut_889_select = {
                             in_data[672],
                             in_data[225],
                             in_data[60],
                             in_data[2],
                             in_data[274],
                             in_data[570]};
    
    wire lut_889_out = lut_889_table[lut_889_select];
    
    generate
    if ( USE_REG ) begin : ff_889
        reg   lut_889_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_889_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_889_ff <= lut_889_out;
            end
        end
        
        assign out_data[889] = lut_889_ff;
    end
    else begin : no_ff_889
        assign out_data[889] = lut_889_out;
    end
    endgenerate
    
    
    
    // LUT : 890
    wire [63:0] lut_890_table = 64'b0000110011001100110001001100110000001100110011001100100011001100;
    wire [5:0] lut_890_select = {
                             in_data[668],
                             in_data[163],
                             in_data[318],
                             in_data[326],
                             in_data[211],
                             in_data[392]};
    
    wire lut_890_out = lut_890_table[lut_890_select];
    
    generate
    if ( USE_REG ) begin : ff_890
        reg   lut_890_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_890_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_890_ff <= lut_890_out;
            end
        end
        
        assign out_data[890] = lut_890_ff;
    end
    else begin : no_ff_890
        assign out_data[890] = lut_890_out;
    end
    endgenerate
    
    
    
    // LUT : 891
    wire [63:0] lut_891_table = 64'b1101110011001111111111001111111111001100110011111100110011001111;
    wire [5:0] lut_891_select = {
                             in_data[704],
                             in_data[110],
                             in_data[495],
                             in_data[633],
                             in_data[260],
                             in_data[448]};
    
    wire lut_891_out = lut_891_table[lut_891_select];
    
    generate
    if ( USE_REG ) begin : ff_891
        reg   lut_891_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_891_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_891_ff <= lut_891_out;
            end
        end
        
        assign out_data[891] = lut_891_ff;
    end
    else begin : no_ff_891
        assign out_data[891] = lut_891_out;
    end
    endgenerate
    
    
    
    // LUT : 892
    wire [63:0] lut_892_table = 64'b0000000000000000000000000000000011111101110111011101110011011100;
    wire [5:0] lut_892_select = {
                             in_data[377],
                             in_data[200],
                             in_data[332],
                             in_data[738],
                             in_data[547],
                             in_data[498]};
    
    wire lut_892_out = lut_892_table[lut_892_select];
    
    generate
    if ( USE_REG ) begin : ff_892
        reg   lut_892_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_892_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_892_ff <= lut_892_out;
            end
        end
        
        assign out_data[892] = lut_892_ff;
    end
    else begin : no_ff_892
        assign out_data[892] = lut_892_out;
    end
    endgenerate
    
    
    
    // LUT : 893
    wire [63:0] lut_893_table = 64'b1111111111111111111111111111111110101110111011101010101010101110;
    wire [5:0] lut_893_select = {
                             in_data[552],
                             in_data[336],
                             in_data[34],
                             in_data[116],
                             in_data[658],
                             in_data[607]};
    
    wire lut_893_out = lut_893_table[lut_893_select];
    
    generate
    if ( USE_REG ) begin : ff_893
        reg   lut_893_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_893_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_893_ff <= lut_893_out;
            end
        end
        
        assign out_data[893] = lut_893_ff;
    end
    else begin : no_ff_893
        assign out_data[893] = lut_893_out;
    end
    endgenerate
    
    
    
    // LUT : 894
    wire [63:0] lut_894_table = 64'b0000000000000000000000000000000001011111010111110101011101010111;
    wire [5:0] lut_894_select = {
                             in_data[346],
                             in_data[172],
                             in_data[420],
                             in_data[574],
                             in_data[700],
                             in_data[740]};
    
    wire lut_894_out = lut_894_table[lut_894_select];
    
    generate
    if ( USE_REG ) begin : ff_894
        reg   lut_894_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_894_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_894_ff <= lut_894_out;
            end
        end
        
        assign out_data[894] = lut_894_ff;
    end
    else begin : no_ff_894
        assign out_data[894] = lut_894_out;
    end
    endgenerate
    
    
    
    // LUT : 895
    wire [63:0] lut_895_table = 64'b1010101011111111101010111111111100000000101000100000000000110010;
    wire [5:0] lut_895_select = {
                             in_data[432],
                             in_data[444],
                             in_data[131],
                             in_data[100],
                             in_data[454],
                             in_data[220]};
    
    wire lut_895_out = lut_895_table[lut_895_select];
    
    generate
    if ( USE_REG ) begin : ff_895
        reg   lut_895_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_895_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_895_ff <= lut_895_out;
            end
        end
        
        assign out_data[895] = lut_895_ff;
    end
    else begin : no_ff_895
        assign out_data[895] = lut_895_out;
    end
    endgenerate
    
    
    
    // LUT : 896
    wire [63:0] lut_896_table = 64'b1011101010101010111110111010101010111010101010101111101010101010;
    wire [5:0] lut_896_select = {
                             in_data[732],
                             in_data[733],
                             in_data[463],
                             in_data[75],
                             in_data[419],
                             in_data[402]};
    
    wire lut_896_out = lut_896_table[lut_896_select];
    
    generate
    if ( USE_REG ) begin : ff_896
        reg   lut_896_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_896_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_896_ff <= lut_896_out;
            end
        end
        
        assign out_data[896] = lut_896_ff;
    end
    else begin : no_ff_896
        assign out_data[896] = lut_896_out;
    end
    endgenerate
    
    
    
    // LUT : 897
    wire [63:0] lut_897_table = 64'b0000000000000000000000000000000001010101010101010101010101010101;
    wire [5:0] lut_897_select = {
                             in_data[333],
                             in_data[12],
                             in_data[481],
                             in_data[88],
                             in_data[617],
                             in_data[604]};
    
    wire lut_897_out = lut_897_table[lut_897_select];
    
    generate
    if ( USE_REG ) begin : ff_897
        reg   lut_897_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_897_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_897_ff <= lut_897_out;
            end
        end
        
        assign out_data[897] = lut_897_ff;
    end
    else begin : no_ff_897
        assign out_data[897] = lut_897_out;
    end
    endgenerate
    
    
    
    // LUT : 898
    wire [63:0] lut_898_table = 64'b1111111100010000111111110001000011110011111100001111001011110000;
    wire [5:0] lut_898_select = {
                             in_data[416],
                             in_data[338],
                             in_data[287],
                             in_data[345],
                             in_data[350],
                             in_data[691]};
    
    wire lut_898_out = lut_898_table[lut_898_select];
    
    generate
    if ( USE_REG ) begin : ff_898
        reg   lut_898_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_898_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_898_ff <= lut_898_out;
            end
        end
        
        assign out_data[898] = lut_898_ff;
    end
    else begin : no_ff_898
        assign out_data[898] = lut_898_out;
    end
    endgenerate
    
    
    
    // LUT : 899
    wire [63:0] lut_899_table = 64'b0000000000000000000000000000010100000000000000000000000000000101;
    wire [5:0] lut_899_select = {
                             in_data[702],
                             in_data[188],
                             in_data[707],
                             in_data[597],
                             in_data[367],
                             in_data[173]};
    
    wire lut_899_out = lut_899_table[lut_899_select];
    
    generate
    if ( USE_REG ) begin : ff_899
        reg   lut_899_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_899_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_899_ff <= lut_899_out;
            end
        end
        
        assign out_data[899] = lut_899_ff;
    end
    else begin : no_ff_899
        assign out_data[899] = lut_899_out;
    end
    endgenerate
    
    
    
    // LUT : 900
    wire [63:0] lut_900_table = 64'b0000000000000000000000000001000100000000000000000000000000010001;
    wire [5:0] lut_900_select = {
                             in_data[5],
                             in_data[496],
                             in_data[122],
                             in_data[558],
                             in_data[566],
                             in_data[536]};
    
    wire lut_900_out = lut_900_table[lut_900_select];
    
    generate
    if ( USE_REG ) begin : ff_900
        reg   lut_900_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_900_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_900_ff <= lut_900_out;
            end
        end
        
        assign out_data[900] = lut_900_ff;
    end
    else begin : no_ff_900
        assign out_data[900] = lut_900_out;
    end
    endgenerate
    
    
    
    // LUT : 901
    wire [63:0] lut_901_table = 64'b0000000000000000001000000010001000000000000000001111001111110010;
    wire [5:0] lut_901_select = {
                             in_data[710],
                             in_data[508],
                             in_data[373],
                             in_data[497],
                             in_data[236],
                             in_data[356]};
    
    wire lut_901_out = lut_901_table[lut_901_select];
    
    generate
    if ( USE_REG ) begin : ff_901
        reg   lut_901_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_901_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_901_ff <= lut_901_out;
            end
        end
        
        assign out_data[901] = lut_901_ff;
    end
    else begin : no_ff_901
        assign out_data[901] = lut_901_out;
    end
    endgenerate
    
    
    
    // LUT : 902
    wire [63:0] lut_902_table = 64'b0000000000000000000000000000000000000001000000110011001100110011;
    wire [5:0] lut_902_select = {
                             in_data[174],
                             in_data[65],
                             in_data[59],
                             in_data[723],
                             in_data[406],
                             in_data[22]};
    
    wire lut_902_out = lut_902_table[lut_902_select];
    
    generate
    if ( USE_REG ) begin : ff_902
        reg   lut_902_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_902_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_902_ff <= lut_902_out;
            end
        end
        
        assign out_data[902] = lut_902_ff;
    end
    else begin : no_ff_902
        assign out_data[902] = lut_902_out;
    end
    endgenerate
    
    
    
    // LUT : 903
    wire [63:0] lut_903_table = 64'b0000000000000000010001000100010001010101000000001101110101000101;
    wire [5:0] lut_903_select = {
                             in_data[299],
                             in_data[337],
                             in_data[696],
                             in_data[224],
                             in_data[47],
                             in_data[362]};
    
    wire lut_903_out = lut_903_table[lut_903_select];
    
    generate
    if ( USE_REG ) begin : ff_903
        reg   lut_903_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_903_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_903_ff <= lut_903_out;
            end
        end
        
        assign out_data[903] = lut_903_ff;
    end
    else begin : no_ff_903
        assign out_data[903] = lut_903_out;
    end
    endgenerate
    
    
    
    // LUT : 904
    wire [63:0] lut_904_table = 64'b1100111111111111000000001000111011001110111111110000000010001110;
    wire [5:0] lut_904_select = {
                             in_data[335],
                             in_data[369],
                             in_data[473],
                             in_data[613],
                             in_data[193],
                             in_data[764]};
    
    wire lut_904_out = lut_904_table[lut_904_select];
    
    generate
    if ( USE_REG ) begin : ff_904
        reg   lut_904_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_904_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_904_ff <= lut_904_out;
            end
        end
        
        assign out_data[904] = lut_904_ff;
    end
    else begin : no_ff_904
        assign out_data[904] = lut_904_out;
    end
    endgenerate
    
    
    
    // LUT : 905
    wire [63:0] lut_905_table = 64'b1111010111110001111100011111001111110011111100111111000111110001;
    wire [5:0] lut_905_select = {
                             in_data[195],
                             in_data[669],
                             in_data[665],
                             in_data[636],
                             in_data[265],
                             in_data[319]};
    
    wire lut_905_out = lut_905_table[lut_905_select];
    
    generate
    if ( USE_REG ) begin : ff_905
        reg   lut_905_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_905_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_905_ff <= lut_905_out;
            end
        end
        
        assign out_data[905] = lut_905_ff;
    end
    else begin : no_ff_905
        assign out_data[905] = lut_905_out;
    end
    endgenerate
    
    
    
    // LUT : 906
    wire [63:0] lut_906_table = 64'b1111111111111111111111111111111111111111111111101111111111111110;
    wire [5:0] lut_906_select = {
                             in_data[453],
                             in_data[645],
                             in_data[446],
                             in_data[471],
                             in_data[534],
                             in_data[50]};
    
    wire lut_906_out = lut_906_table[lut_906_select];
    
    generate
    if ( USE_REG ) begin : ff_906
        reg   lut_906_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_906_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_906_ff <= lut_906_out;
            end
        end
        
        assign out_data[906] = lut_906_ff;
    end
    else begin : no_ff_906
        assign out_data[906] = lut_906_out;
    end
    endgenerate
    
    
    
    // LUT : 907
    wire [63:0] lut_907_table = 64'b1011101110111011111110101011101010111011101110111011101010111010;
    wire [5:0] lut_907_select = {
                             in_data[73],
                             in_data[320],
                             in_data[61],
                             in_data[395],
                             in_data[708],
                             in_data[405]};
    
    wire lut_907_out = lut_907_table[lut_907_select];
    
    generate
    if ( USE_REG ) begin : ff_907
        reg   lut_907_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_907_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_907_ff <= lut_907_out;
            end
        end
        
        assign out_data[907] = lut_907_ff;
    end
    else begin : no_ff_907
        assign out_data[907] = lut_907_out;
    end
    endgenerate
    
    
    
    // LUT : 908
    wire [63:0] lut_908_table = 64'b0000000000000000111111111111111100000000000000001111111111111111;
    wire [5:0] lut_908_select = {
                             in_data[701],
                             in_data[515],
                             in_data[624],
                             in_data[58],
                             in_data[83],
                             in_data[151]};
    
    wire lut_908_out = lut_908_table[lut_908_select];
    
    generate
    if ( USE_REG ) begin : ff_908
        reg   lut_908_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_908_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_908_ff <= lut_908_out;
            end
        end
        
        assign out_data[908] = lut_908_ff;
    end
    else begin : no_ff_908
        assign out_data[908] = lut_908_out;
    end
    endgenerate
    
    
    
    // LUT : 909
    wire [63:0] lut_909_table = 64'b0001010101010101000001010000010100010101000101010000010100000101;
    wire [5:0] lut_909_select = {
                             in_data[538],
                             in_data[44],
                             in_data[729],
                             in_data[330],
                             in_data[366],
                             in_data[690]};
    
    wire lut_909_out = lut_909_table[lut_909_select];
    
    generate
    if ( USE_REG ) begin : ff_909
        reg   lut_909_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_909_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_909_ff <= lut_909_out;
            end
        end
        
        assign out_data[909] = lut_909_ff;
    end
    else begin : no_ff_909
        assign out_data[909] = lut_909_out;
    end
    endgenerate
    
    
    
    // LUT : 910
    wire [63:0] lut_910_table = 64'b0000000100000001000000010000000100000111000001110001001100010011;
    wire [5:0] lut_910_select = {
                             in_data[119],
                             in_data[383],
                             in_data[143],
                             in_data[465],
                             in_data[389],
                             in_data[118]};
    
    wire lut_910_out = lut_910_table[lut_910_select];
    
    generate
    if ( USE_REG ) begin : ff_910
        reg   lut_910_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_910_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_910_ff <= lut_910_out;
            end
        end
        
        assign out_data[910] = lut_910_ff;
    end
    else begin : no_ff_910
        assign out_data[910] = lut_910_out;
    end
    endgenerate
    
    
    
    // LUT : 911
    wire [63:0] lut_911_table = 64'b0000000000001111000000000000000100000000111111110000000011111111;
    wire [5:0] lut_911_select = {
                             in_data[571],
                             in_data[152],
                             in_data[490],
                             in_data[477],
                             in_data[599],
                             in_data[754]};
    
    wire lut_911_out = lut_911_table[lut_911_select];
    
    generate
    if ( USE_REG ) begin : ff_911
        reg   lut_911_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_911_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_911_ff <= lut_911_out;
            end
        end
        
        assign out_data[911] = lut_911_ff;
    end
    else begin : no_ff_911
        assign out_data[911] = lut_911_out;
    end
    endgenerate
    
    
    
    // LUT : 912
    wire [63:0] lut_912_table = 64'b1111111111111111000000000000000011110000111111110000000011111111;
    wire [5:0] lut_912_select = {
                             in_data[429],
                             in_data[694],
                             in_data[398],
                             in_data[377],
                             in_data[43],
                             in_data[586]};
    
    wire lut_912_out = lut_912_table[lut_912_select];
    
    generate
    if ( USE_REG ) begin : ff_912
        reg   lut_912_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_912_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_912_ff <= lut_912_out;
            end
        end
        
        assign out_data[912] = lut_912_ff;
    end
    else begin : no_ff_912
        assign out_data[912] = lut_912_out;
    end
    endgenerate
    
    
    
    // LUT : 913
    wire [63:0] lut_913_table = 64'b0101010101010101111111110101010101010101010101010101010101010101;
    wire [5:0] lut_913_select = {
                             in_data[67],
                             in_data[581],
                             in_data[716],
                             in_data[764],
                             in_data[86],
                             in_data[216]};
    
    wire lut_913_out = lut_913_table[lut_913_select];
    
    generate
    if ( USE_REG ) begin : ff_913
        reg   lut_913_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_913_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_913_ff <= lut_913_out;
            end
        end
        
        assign out_data[913] = lut_913_ff;
    end
    else begin : no_ff_913
        assign out_data[913] = lut_913_out;
    end
    endgenerate
    
    
    
    // LUT : 914
    wire [63:0] lut_914_table = 64'b1111111111111111000000000000000011111111111111110100010001001100;
    wire [5:0] lut_914_select = {
                             in_data[706],
                             in_data[664],
                             in_data[592],
                             in_data[54],
                             in_data[558],
                             in_data[507]};
    
    wire lut_914_out = lut_914_table[lut_914_select];
    
    generate
    if ( USE_REG ) begin : ff_914
        reg   lut_914_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_914_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_914_ff <= lut_914_out;
            end
        end
        
        assign out_data[914] = lut_914_ff;
    end
    else begin : no_ff_914
        assign out_data[914] = lut_914_out;
    end
    endgenerate
    
    
    
    // LUT : 915
    wire [63:0] lut_915_table = 64'b1110110011111110110011001111110011111100111111111111110011111110;
    wire [5:0] lut_915_select = {
                             in_data[193],
                             in_data[76],
                             in_data[608],
                             in_data[302],
                             in_data[122],
                             in_data[451]};
    
    wire lut_915_out = lut_915_table[lut_915_select];
    
    generate
    if ( USE_REG ) begin : ff_915
        reg   lut_915_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_915_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_915_ff <= lut_915_out;
            end
        end
        
        assign out_data[915] = lut_915_ff;
    end
    else begin : no_ff_915
        assign out_data[915] = lut_915_out;
    end
    endgenerate
    
    
    
    // LUT : 916
    wire [63:0] lut_916_table = 64'b0100010100000101000001010000000011110101111101011111010111110101;
    wire [5:0] lut_916_select = {
                             in_data[425],
                             in_data[26],
                             in_data[501],
                             in_data[205],
                             in_data[336],
                             in_data[357]};
    
    wire lut_916_out = lut_916_table[lut_916_select];
    
    generate
    if ( USE_REG ) begin : ff_916
        reg   lut_916_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_916_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_916_ff <= lut_916_out;
            end
        end
        
        assign out_data[916] = lut_916_ff;
    end
    else begin : no_ff_916
        assign out_data[916] = lut_916_out;
    end
    endgenerate
    
    
    
    // LUT : 917
    wire [63:0] lut_917_table = 64'b1111111111111101111111111101110111111111110011001111110111011100;
    wire [5:0] lut_917_select = {
                             in_data[483],
                             in_data[346],
                             in_data[153],
                             in_data[63],
                             in_data[330],
                             in_data[433]};
    
    wire lut_917_out = lut_917_table[lut_917_select];
    
    generate
    if ( USE_REG ) begin : ff_917
        reg   lut_917_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_917_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_917_ff <= lut_917_out;
            end
        end
        
        assign out_data[917] = lut_917_ff;
    end
    else begin : no_ff_917
        assign out_data[917] = lut_917_out;
    end
    endgenerate
    
    
    
    // LUT : 918
    wire [63:0] lut_918_table = 64'b0000111100000000000011110000000011111111000011001100111100001100;
    wire [5:0] lut_918_select = {
                             in_data[709],
                             in_data[280],
                             in_data[566],
                             in_data[715],
                             in_data[222],
                             in_data[141]};
    
    wire lut_918_out = lut_918_table[lut_918_select];
    
    generate
    if ( USE_REG ) begin : ff_918
        reg   lut_918_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_918_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_918_ff <= lut_918_out;
            end
        end
        
        assign out_data[918] = lut_918_ff;
    end
    else begin : no_ff_918
        assign out_data[918] = lut_918_out;
    end
    endgenerate
    
    
    
    // LUT : 919
    wire [63:0] lut_919_table = 64'b1111111101010000111111010000000011111111010101001111010101010000;
    wire [5:0] lut_919_select = {
                             in_data[130],
                             in_data[172],
                             in_data[375],
                             in_data[278],
                             in_data[40],
                             in_data[611]};
    
    wire lut_919_out = lut_919_table[lut_919_select];
    
    generate
    if ( USE_REG ) begin : ff_919
        reg   lut_919_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_919_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_919_ff <= lut_919_out;
            end
        end
        
        assign out_data[919] = lut_919_ff;
    end
    else begin : no_ff_919
        assign out_data[919] = lut_919_out;
    end
    endgenerate
    
    
    
    // LUT : 920
    wire [63:0] lut_920_table = 64'b1101010111010100111111011111110111010100110101001111110111111101;
    wire [5:0] lut_920_select = {
                             in_data[618],
                             in_data[292],
                             in_data[755],
                             in_data[583],
                             in_data[369],
                             in_data[604]};
    
    wire lut_920_out = lut_920_table[lut_920_select];
    
    generate
    if ( USE_REG ) begin : ff_920
        reg   lut_920_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_920_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_920_ff <= lut_920_out;
            end
        end
        
        assign out_data[920] = lut_920_ff;
    end
    else begin : no_ff_920
        assign out_data[920] = lut_920_out;
    end
    endgenerate
    
    
    
    // LUT : 921
    wire [63:0] lut_921_table = 64'b1111000011110001000000000000000011110000111100010000000000000000;
    wire [5:0] lut_921_select = {
                             in_data[531],
                             in_data[352],
                             in_data[394],
                             in_data[349],
                             in_data[609],
                             in_data[728]};
    
    wire lut_921_out = lut_921_table[lut_921_select];
    
    generate
    if ( USE_REG ) begin : ff_921
        reg   lut_921_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_921_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_921_ff <= lut_921_out;
            end
        end
        
        assign out_data[921] = lut_921_ff;
    end
    else begin : no_ff_921
        assign out_data[921] = lut_921_out;
    end
    endgenerate
    
    
    
    // LUT : 922
    wire [63:0] lut_922_table = 64'b1111111111111111111100001111000011111111111111111111000011110000;
    wire [5:0] lut_922_select = {
                             in_data[17],
                             in_data[712],
                             in_data[475],
                             in_data[347],
                             in_data[89],
                             in_data[70]};
    
    wire lut_922_out = lut_922_table[lut_922_select];
    
    generate
    if ( USE_REG ) begin : ff_922
        reg   lut_922_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_922_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_922_ff <= lut_922_out;
            end
        end
        
        assign out_data[922] = lut_922_ff;
    end
    else begin : no_ff_922
        assign out_data[922] = lut_922_out;
    end
    endgenerate
    
    
    
    // LUT : 923
    wire [63:0] lut_923_table = 64'b0000000000100000000000000001000011110000111100001111000011110000;
    wire [5:0] lut_923_select = {
                             in_data[550],
                             in_data[700],
                             in_data[750],
                             in_data[214],
                             in_data[773],
                             in_data[27]};
    
    wire lut_923_out = lut_923_table[lut_923_select];
    
    generate
    if ( USE_REG ) begin : ff_923
        reg   lut_923_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_923_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_923_ff <= lut_923_out;
            end
        end
        
        assign out_data[923] = lut_923_ff;
    end
    else begin : no_ff_923
        assign out_data[923] = lut_923_out;
    end
    endgenerate
    
    
    
    // LUT : 924
    wire [63:0] lut_924_table = 64'b0100010000000000111011101010101001000100000000001110111010101010;
    wire [5:0] lut_924_select = {
                             in_data[617],
                             in_data[179],
                             in_data[406],
                             in_data[530],
                             in_data[331],
                             in_data[326]};
    
    wire lut_924_out = lut_924_table[lut_924_select];
    
    generate
    if ( USE_REG ) begin : ff_924
        reg   lut_924_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_924_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_924_ff <= lut_924_out;
            end
        end
        
        assign out_data[924] = lut_924_ff;
    end
    else begin : no_ff_924
        assign out_data[924] = lut_924_out;
    end
    endgenerate
    
    
    
    // LUT : 925
    wire [63:0] lut_925_table = 64'b1100000011000000111000001100000011100000111000001111000011100000;
    wire [5:0] lut_925_select = {
                             in_data[536],
                             in_data[38],
                             in_data[224],
                             in_data[461],
                             in_data[460],
                             in_data[195]};
    
    wire lut_925_out = lut_925_table[lut_925_select];
    
    generate
    if ( USE_REG ) begin : ff_925
        reg   lut_925_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_925_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_925_ff <= lut_925_out;
            end
        end
        
        assign out_data[925] = lut_925_ff;
    end
    else begin : no_ff_925
        assign out_data[925] = lut_925_out;
    end
    endgenerate
    
    
    
    // LUT : 926
    wire [63:0] lut_926_table = 64'b0000000001011111000000000111111100000000111100000000000011110000;
    wire [5:0] lut_926_select = {
                             in_data[509],
                             in_data[420],
                             in_data[177],
                             in_data[484],
                             in_data[225],
                             in_data[693]};
    
    wire lut_926_out = lut_926_table[lut_926_select];
    
    generate
    if ( USE_REG ) begin : ff_926
        reg   lut_926_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_926_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_926_ff <= lut_926_out;
            end
        end
        
        assign out_data[926] = lut_926_ff;
    end
    else begin : no_ff_926
        assign out_data[926] = lut_926_out;
    end
    endgenerate
    
    
    
    // LUT : 927
    wire [63:0] lut_927_table = 64'b1110111011001100111011101000110011111111111011101111111111101111;
    wire [5:0] lut_927_select = {
                             in_data[680],
                             in_data[11],
                             in_data[229],
                             in_data[668],
                             in_data[50],
                             in_data[64]};
    
    wire lut_927_out = lut_927_table[lut_927_select];
    
    generate
    if ( USE_REG ) begin : ff_927
        reg   lut_927_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_927_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_927_ff <= lut_927_out;
            end
        end
        
        assign out_data[927] = lut_927_ff;
    end
    else begin : no_ff_927
        assign out_data[927] = lut_927_out;
    end
    endgenerate
    
    
    
    // LUT : 928
    wire [63:0] lut_928_table = 64'b0000000000000010000000000000000000000011001000110000000100011111;
    wire [5:0] lut_928_select = {
                             in_data[206],
                             in_data[370],
                             in_data[707],
                             in_data[691],
                             in_data[714],
                             in_data[576]};
    
    wire lut_928_out = lut_928_table[lut_928_select];
    
    generate
    if ( USE_REG ) begin : ff_928
        reg   lut_928_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_928_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_928_ff <= lut_928_out;
            end
        end
        
        assign out_data[928] = lut_928_ff;
    end
    else begin : no_ff_928
        assign out_data[928] = lut_928_out;
    end
    endgenerate
    
    
    
    // LUT : 929
    wire [63:0] lut_929_table = 64'b1111010011110100111101011111010100000000000000000001000100110001;
    wire [5:0] lut_929_select = {
                             in_data[434],
                             in_data[685],
                             in_data[758],
                             in_data[293],
                             in_data[316],
                             in_data[464]};
    
    wire lut_929_out = lut_929_table[lut_929_select];
    
    generate
    if ( USE_REG ) begin : ff_929
        reg   lut_929_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_929_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_929_ff <= lut_929_out;
            end
        end
        
        assign out_data[929] = lut_929_ff;
    end
    else begin : no_ff_929
        assign out_data[929] = lut_929_out;
    end
    endgenerate
    
    
    
    // LUT : 930
    wire [63:0] lut_930_table = 64'b0000000100000000000000010000000000010011000100110001001100010011;
    wire [5:0] lut_930_select = {
                             in_data[512],
                             in_data[84],
                             in_data[323],
                             in_data[546],
                             in_data[516],
                             in_data[81]};
    
    wire lut_930_out = lut_930_table[lut_930_select];
    
    generate
    if ( USE_REG ) begin : ff_930
        reg   lut_930_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_930_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_930_ff <= lut_930_out;
            end
        end
        
        assign out_data[930] = lut_930_ff;
    end
    else begin : no_ff_930
        assign out_data[930] = lut_930_out;
    end
    endgenerate
    
    
    
    // LUT : 931
    wire [63:0] lut_931_table = 64'b1111111111111111111111111111111111111111111011110000000000000000;
    wire [5:0] lut_931_select = {
                             in_data[564],
                             in_data[208],
                             in_data[178],
                             in_data[47],
                             in_data[129],
                             in_data[80]};
    
    wire lut_931_out = lut_931_table[lut_931_select];
    
    generate
    if ( USE_REG ) begin : ff_931
        reg   lut_931_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_931_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_931_ff <= lut_931_out;
            end
        end
        
        assign out_data[931] = lut_931_ff;
    end
    else begin : no_ff_931
        assign out_data[931] = lut_931_out;
    end
    endgenerate
    
    
    
    // LUT : 932
    wire [63:0] lut_932_table = 64'b1000100010001000111011101110111000000000000000001111111011111110;
    wire [5:0] lut_932_select = {
                             in_data[159],
                             in_data[652],
                             in_data[110],
                             in_data[743],
                             in_data[97],
                             in_data[413]};
    
    wire lut_932_out = lut_932_table[lut_932_select];
    
    generate
    if ( USE_REG ) begin : ff_932
        reg   lut_932_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_932_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_932_ff <= lut_932_out;
            end
        end
        
        assign out_data[932] = lut_932_ff;
    end
    else begin : no_ff_932
        assign out_data[932] = lut_932_out;
    end
    endgenerate
    
    
    
    // LUT : 933
    wire [63:0] lut_933_table = 64'b0000000001000100000000000100010000000000110111010000000011011101;
    wire [5:0] lut_933_select = {
                             in_data[747],
                             in_data[757],
                             in_data[416],
                             in_data[21],
                             in_data[527],
                             in_data[543]};
    
    wire lut_933_out = lut_933_table[lut_933_select];
    
    generate
    if ( USE_REG ) begin : ff_933
        reg   lut_933_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_933_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_933_ff <= lut_933_out;
            end
        end
        
        assign out_data[933] = lut_933_ff;
    end
    else begin : no_ff_933
        assign out_data[933] = lut_933_out;
    end
    endgenerate
    
    
    
    // LUT : 934
    wire [63:0] lut_934_table = 64'b1111111111111111111111100000110011111111111111111111111100001100;
    wire [5:0] lut_934_select = {
                             in_data[22],
                             in_data[262],
                             in_data[596],
                             in_data[468],
                             in_data[740],
                             in_data[724]};
    
    wire lut_934_out = lut_934_table[lut_934_select];
    
    generate
    if ( USE_REG ) begin : ff_934
        reg   lut_934_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_934_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_934_ff <= lut_934_out;
            end
        end
        
        assign out_data[934] = lut_934_ff;
    end
    else begin : no_ff_934
        assign out_data[934] = lut_934_out;
    end
    endgenerate
    
    
    
    // LUT : 935
    wire [63:0] lut_935_table = 64'b0000000000000000011100010111000100000000000000000111000101110001;
    wire [5:0] lut_935_select = {
                             in_data[82],
                             in_data[244],
                             in_data[616],
                             in_data[339],
                             in_data[414],
                             in_data[649]};
    
    wire lut_935_out = lut_935_table[lut_935_select];
    
    generate
    if ( USE_REG ) begin : ff_935
        reg   lut_935_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_935_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_935_ff <= lut_935_out;
            end
        end
        
        assign out_data[935] = lut_935_ff;
    end
    else begin : no_ff_935
        assign out_data[935] = lut_935_out;
    end
    endgenerate
    
    
    
    // LUT : 936
    wire [63:0] lut_936_table = 64'b0000000000000000000000000000000000000000000000001111011111111111;
    wire [5:0] lut_936_select = {
                             in_data[215],
                             in_data[299],
                             in_data[335],
                             in_data[761],
                             in_data[573],
                             in_data[521]};
    
    wire lut_936_out = lut_936_table[lut_936_select];
    
    generate
    if ( USE_REG ) begin : ff_936
        reg   lut_936_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_936_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_936_ff <= lut_936_out;
            end
        end
        
        assign out_data[936] = lut_936_ff;
    end
    else begin : no_ff_936
        assign out_data[936] = lut_936_out;
    end
    endgenerate
    
    
    
    // LUT : 937
    wire [63:0] lut_937_table = 64'b0101010101000101010101010101010101010101000000001111111101010101;
    wire [5:0] lut_937_select = {
                             in_data[241],
                             in_data[582],
                             in_data[517],
                             in_data[478],
                             in_data[600],
                             in_data[212]};
    
    wire lut_937_out = lut_937_table[lut_937_select];
    
    generate
    if ( USE_REG ) begin : ff_937
        reg   lut_937_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_937_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_937_ff <= lut_937_out;
            end
        end
        
        assign out_data[937] = lut_937_ff;
    end
    else begin : no_ff_937
        assign out_data[937] = lut_937_out;
    end
    endgenerate
    
    
    
    // LUT : 938
    wire [63:0] lut_938_table = 64'b0000000000001010000000001010111100000000000011110000000000101111;
    wire [5:0] lut_938_select = {
                             in_data[471],
                             in_data[271],
                             in_data[480],
                             in_data[486],
                             in_data[113],
                             in_data[145]};
    
    wire lut_938_out = lut_938_table[lut_938_select];
    
    generate
    if ( USE_REG ) begin : ff_938
        reg   lut_938_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_938_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_938_ff <= lut_938_out;
            end
        end
        
        assign out_data[938] = lut_938_ff;
    end
    else begin : no_ff_938
        assign out_data[938] = lut_938_out;
    end
    endgenerate
    
    
    
    // LUT : 939
    wire [63:0] lut_939_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_939_select = {
                             in_data[197],
                             in_data[380],
                             in_data[771],
                             in_data[458],
                             in_data[646],
                             in_data[16]};
    
    wire lut_939_out = lut_939_table[lut_939_select];
    
    generate
    if ( USE_REG ) begin : ff_939
        reg   lut_939_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_939_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_939_ff <= lut_939_out;
            end
        end
        
        assign out_data[939] = lut_939_ff;
    end
    else begin : no_ff_939
        assign out_data[939] = lut_939_out;
    end
    endgenerate
    
    
    
    // LUT : 940
    wire [63:0] lut_940_table = 64'b0000000011111111000000000111011100000000111111110000000011111111;
    wire [5:0] lut_940_select = {
                             in_data[114],
                             in_data[588],
                             in_data[345],
                             in_data[777],
                             in_data[597],
                             in_data[137]};
    
    wire lut_940_out = lut_940_table[lut_940_select];
    
    generate
    if ( USE_REG ) begin : ff_940
        reg   lut_940_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_940_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_940_ff <= lut_940_out;
            end
        end
        
        assign out_data[940] = lut_940_ff;
    end
    else begin : no_ff_940
        assign out_data[940] = lut_940_out;
    end
    endgenerate
    
    
    
    // LUT : 941
    wire [63:0] lut_941_table = 64'b0000000000000000111111111111111100000000110011001111111111111111;
    wire [5:0] lut_941_select = {
                             in_data[628],
                             in_data[542],
                             in_data[147],
                             in_data[447],
                             in_data[631],
                             in_data[228]};
    
    wire lut_941_out = lut_941_table[lut_941_select];
    
    generate
    if ( USE_REG ) begin : ff_941
        reg   lut_941_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_941_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_941_ff <= lut_941_out;
            end
        end
        
        assign out_data[941] = lut_941_ff;
    end
    else begin : no_ff_941
        assign out_data[941] = lut_941_out;
    end
    endgenerate
    
    
    
    // LUT : 942
    wire [63:0] lut_942_table = 64'b1000111011111111000010000000111010101111111111110000100000001110;
    wire [5:0] lut_942_select = {
                             in_data[73],
                             in_data[683],
                             in_data[259],
                             in_data[312],
                             in_data[117],
                             in_data[630]};
    
    wire lut_942_out = lut_942_table[lut_942_select];
    
    generate
    if ( USE_REG ) begin : ff_942
        reg   lut_942_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_942_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_942_ff <= lut_942_out;
            end
        end
        
        assign out_data[942] = lut_942_ff;
    end
    else begin : no_ff_942
        assign out_data[942] = lut_942_out;
    end
    endgenerate
    
    
    
    // LUT : 943
    wire [63:0] lut_943_table = 64'b1010101111111011101010101010101011111111101010101010101010101010;
    wire [5:0] lut_943_select = {
                             in_data[538],
                             in_data[282],
                             in_data[182],
                             in_data[340],
                             in_data[696],
                             in_data[602]};
    
    wire lut_943_out = lut_943_table[lut_943_select];
    
    generate
    if ( USE_REG ) begin : ff_943
        reg   lut_943_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_943_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_943_ff <= lut_943_out;
            end
        end
        
        assign out_data[943] = lut_943_ff;
    end
    else begin : no_ff_943
        assign out_data[943] = lut_943_out;
    end
    endgenerate
    
    
    
    // LUT : 944
    wire [63:0] lut_944_table = 64'b0000000000000000000000000000010100000000000000000000000000000111;
    wire [5:0] lut_944_select = {
                             in_data[171],
                             in_data[635],
                             in_data[595],
                             in_data[660],
                             in_data[614],
                             in_data[92]};
    
    wire lut_944_out = lut_944_table[lut_944_select];
    
    generate
    if ( USE_REG ) begin : ff_944
        reg   lut_944_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_944_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_944_ff <= lut_944_out;
            end
        end
        
        assign out_data[944] = lut_944_ff;
    end
    else begin : no_ff_944
        assign out_data[944] = lut_944_out;
    end
    endgenerate
    
    
    
    // LUT : 945
    wire [63:0] lut_945_table = 64'b1111111111111111000000001100111111111111111111110000000000000000;
    wire [5:0] lut_945_select = {
                             in_data[513],
                             in_data[496],
                             in_data[237],
                             in_data[277],
                             in_data[18],
                             in_data[7]};
    
    wire lut_945_out = lut_945_table[lut_945_select];
    
    generate
    if ( USE_REG ) begin : ff_945
        reg   lut_945_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_945_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_945_ff <= lut_945_out;
            end
        end
        
        assign out_data[945] = lut_945_ff;
    end
    else begin : no_ff_945
        assign out_data[945] = lut_945_out;
    end
    endgenerate
    
    
    
    // LUT : 946
    wire [63:0] lut_946_table = 64'b0000000000000100010001001100110011011100110011001111111111001100;
    wire [5:0] lut_946_select = {
                             in_data[128],
                             in_data[367],
                             in_data[372],
                             in_data[734],
                             in_data[246],
                             in_data[65]};
    
    wire lut_946_out = lut_946_table[lut_946_select];
    
    generate
    if ( USE_REG ) begin : ff_946
        reg   lut_946_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_946_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_946_ff <= lut_946_out;
            end
        end
        
        assign out_data[946] = lut_946_ff;
    end
    else begin : no_ff_946
        assign out_data[946] = lut_946_out;
    end
    endgenerate
    
    
    
    // LUT : 947
    wire [63:0] lut_947_table = 64'b0000000000000000000000000000000000000001000000010000000100000011;
    wire [5:0] lut_947_select = {
                             in_data[120],
                             in_data[167],
                             in_data[165],
                             in_data[637],
                             in_data[624],
                             in_data[258]};
    
    wire lut_947_out = lut_947_table[lut_947_select];
    
    generate
    if ( USE_REG ) begin : ff_947
        reg   lut_947_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_947_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_947_ff <= lut_947_out;
            end
        end
        
        assign out_data[947] = lut_947_ff;
    end
    else begin : no_ff_947
        assign out_data[947] = lut_947_out;
    end
    endgenerate
    
    
    
    // LUT : 948
    wire [63:0] lut_948_table = 64'b0000000000000000000000000000000000000101000001010000010100000101;
    wire [5:0] lut_948_select = {
                             in_data[180],
                             in_data[226],
                             in_data[421],
                             in_data[284],
                             in_data[33],
                             in_data[679]};
    
    wire lut_948_out = lut_948_table[lut_948_select];
    
    generate
    if ( USE_REG ) begin : ff_948
        reg   lut_948_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_948_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_948_ff <= lut_948_out;
            end
        end
        
        assign out_data[948] = lut_948_ff;
    end
    else begin : no_ff_948
        assign out_data[948] = lut_948_out;
    end
    endgenerate
    
    
    
    // LUT : 949
    wire [63:0] lut_949_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_949_select = {
                             in_data[391],
                             in_data[88],
                             in_data[762],
                             in_data[674],
                             in_data[437],
                             in_data[540]};
    
    wire lut_949_out = lut_949_table[lut_949_select];
    
    generate
    if ( USE_REG ) begin : ff_949
        reg   lut_949_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_949_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_949_ff <= lut_949_out;
            end
        end
        
        assign out_data[949] = lut_949_ff;
    end
    else begin : no_ff_949
        assign out_data[949] = lut_949_out;
    end
    endgenerate
    
    
    
    // LUT : 950
    wire [63:0] lut_950_table = 64'b1111111111111111111111101111111111111111111111111111111011111110;
    wire [5:0] lut_950_select = {
                             in_data[502],
                             in_data[650],
                             in_data[725],
                             in_data[470],
                             in_data[622],
                             in_data[102]};
    
    wire lut_950_out = lut_950_table[lut_950_select];
    
    generate
    if ( USE_REG ) begin : ff_950
        reg   lut_950_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_950_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_950_ff <= lut_950_out;
            end
        end
        
        assign out_data[950] = lut_950_ff;
    end
    else begin : no_ff_950
        assign out_data[950] = lut_950_out;
    end
    endgenerate
    
    
    
    // LUT : 951
    wire [63:0] lut_951_table = 64'b0000000000001010000000000000101100001010000010100000001000001111;
    wire [5:0] lut_951_select = {
                             in_data[68],
                             in_data[231],
                             in_data[711],
                             in_data[654],
                             in_data[473],
                             in_data[663]};
    
    wire lut_951_out = lut_951_table[lut_951_select];
    
    generate
    if ( USE_REG ) begin : ff_951
        reg   lut_951_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_951_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_951_ff <= lut_951_out;
            end
        end
        
        assign out_data[951] = lut_951_ff;
    end
    else begin : no_ff_951
        assign out_data[951] = lut_951_out;
    end
    endgenerate
    
    
    
    // LUT : 952
    wire [63:0] lut_952_table = 64'b1100000011100000110011101111111111001000111000001100111011111111;
    wire [5:0] lut_952_select = {
                             in_data[71],
                             in_data[603],
                             in_data[234],
                             in_data[121],
                             in_data[488],
                             in_data[390]};
    
    wire lut_952_out = lut_952_table[lut_952_select];
    
    generate
    if ( USE_REG ) begin : ff_952
        reg   lut_952_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_952_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_952_ff <= lut_952_out;
            end
        end
        
        assign out_data[952] = lut_952_ff;
    end
    else begin : no_ff_952
        assign out_data[952] = lut_952_out;
    end
    endgenerate
    
    
    
    // LUT : 953
    wire [63:0] lut_953_table = 64'b1111000011110011111100001111001111110000111100111111000011110011;
    wire [5:0] lut_953_select = {
                             in_data[642],
                             in_data[45],
                             in_data[242],
                             in_data[360],
                             in_data[733],
                             in_data[79]};
    
    wire lut_953_out = lut_953_table[lut_953_select];
    
    generate
    if ( USE_REG ) begin : ff_953
        reg   lut_953_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_953_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_953_ff <= lut_953_out;
            end
        end
        
        assign out_data[953] = lut_953_ff;
    end
    else begin : no_ff_953
        assign out_data[953] = lut_953_out;
    end
    endgenerate
    
    
    
    // LUT : 954
    wire [63:0] lut_954_table = 64'b0111011101110110011101110111011001110101011101100111011101110110;
    wire [5:0] lut_954_select = {
                             in_data[708],
                             in_data[769],
                             in_data[522],
                             in_data[499],
                             in_data[511],
                             in_data[457]};
    
    wire lut_954_out = lut_954_table[lut_954_select];
    
    generate
    if ( USE_REG ) begin : ff_954
        reg   lut_954_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_954_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_954_ff <= lut_954_out;
            end
        end
        
        assign out_data[954] = lut_954_ff;
    end
    else begin : no_ff_954
        assign out_data[954] = lut_954_out;
    end
    endgenerate
    
    
    
    // LUT : 955
    wire [63:0] lut_955_table = 64'b1010111010101110111011101110111010101010101010101110111011101110;
    wire [5:0] lut_955_select = {
                             in_data[199],
                             in_data[395],
                             in_data[767],
                             in_data[55],
                             in_data[574],
                             in_data[127]};
    
    wire lut_955_out = lut_955_table[lut_955_select];
    
    generate
    if ( USE_REG ) begin : ff_955
        reg   lut_955_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_955_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_955_ff <= lut_955_out;
            end
        end
        
        assign out_data[955] = lut_955_ff;
    end
    else begin : no_ff_955
        assign out_data[955] = lut_955_out;
    end
    endgenerate
    
    
    
    // LUT : 956
    wire [63:0] lut_956_table = 64'b0000000011111111111110001111100010100000111111111111101011111111;
    wire [5:0] lut_956_select = {
                             in_data[446],
                             in_data[131],
                             in_data[657],
                             in_data[396],
                             in_data[78],
                             in_data[90]};
    
    wire lut_956_out = lut_956_table[lut_956_select];
    
    generate
    if ( USE_REG ) begin : ff_956
        reg   lut_956_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_956_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_956_ff <= lut_956_out;
            end
        end
        
        assign out_data[956] = lut_956_ff;
    end
    else begin : no_ff_956
        assign out_data[956] = lut_956_out;
    end
    endgenerate
    
    
    
    // LUT : 957
    wire [63:0] lut_957_table = 64'b1111111110111111111111110010111111111111101111111111111100101111;
    wire [5:0] lut_957_select = {
                             in_data[772],
                             in_data[658],
                             in_data[686],
                             in_data[489],
                             in_data[621],
                             in_data[104]};
    
    wire lut_957_out = lut_957_table[lut_957_select];
    
    generate
    if ( USE_REG ) begin : ff_957
        reg   lut_957_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_957_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_957_ff <= lut_957_out;
            end
        end
        
        assign out_data[957] = lut_957_ff;
    end
    else begin : no_ff_957
        assign out_data[957] = lut_957_out;
    end
    endgenerate
    
    
    
    // LUT : 958
    wire [63:0] lut_958_table = 64'b0000000000000000000100010001001100000000000000000001000100010011;
    wire [5:0] lut_958_select = {
                             in_data[9],
                             in_data[682],
                             in_data[452],
                             in_data[426],
                             in_data[238],
                             in_data[322]};
    
    wire lut_958_out = lut_958_table[lut_958_select];
    
    generate
    if ( USE_REG ) begin : ff_958
        reg   lut_958_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_958_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_958_ff <= lut_958_out;
            end
        end
        
        assign out_data[958] = lut_958_ff;
    end
    else begin : no_ff_958
        assign out_data[958] = lut_958_out;
    end
    endgenerate
    
    
    
    // LUT : 959
    wire [63:0] lut_959_table = 64'b0111000011110000101000001111000011111010111110101111101011111010;
    wire [5:0] lut_959_select = {
                             in_data[405],
                             in_data[569],
                             in_data[3],
                             in_data[577],
                             in_data[732],
                             in_data[155]};
    
    wire lut_959_out = lut_959_table[lut_959_select];
    
    generate
    if ( USE_REG ) begin : ff_959
        reg   lut_959_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_959_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_959_ff <= lut_959_out;
            end
        end
        
        assign out_data[959] = lut_959_ff;
    end
    else begin : no_ff_959
        assign out_data[959] = lut_959_out;
    end
    endgenerate
    
    
    
    // LUT : 960
    wire [63:0] lut_960_table = 64'b0011111100000000001100110000000011111111011101111111111100110011;
    wire [5:0] lut_960_select = {
                             in_data[350],
                             in_data[173],
                             in_data[387],
                             in_data[297],
                             in_data[181],
                             in_data[106]};
    
    wire lut_960_out = lut_960_table[lut_960_select];
    
    generate
    if ( USE_REG ) begin : ff_960
        reg   lut_960_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_960_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_960_ff <= lut_960_out;
            end
        end
        
        assign out_data[960] = lut_960_ff;
    end
    else begin : no_ff_960
        assign out_data[960] = lut_960_out;
    end
    endgenerate
    
    
    
    // LUT : 961
    wire [63:0] lut_961_table = 64'b1111111111111111111111111111111111111111111111110000000011010100;
    wire [5:0] lut_961_select = {
                             in_data[93],
                             in_data[626],
                             in_data[427],
                             in_data[28],
                             in_data[697],
                             in_data[373]};
    
    wire lut_961_out = lut_961_table[lut_961_select];
    
    generate
    if ( USE_REG ) begin : ff_961
        reg   lut_961_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_961_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_961_ff <= lut_961_out;
            end
        end
        
        assign out_data[961] = lut_961_ff;
    end
    else begin : no_ff_961
        assign out_data[961] = lut_961_out;
    end
    endgenerate
    
    
    
    // LUT : 962
    wire [63:0] lut_962_table = 64'b1100111100001111110011110000111111001111000011001100111100001111;
    wire [5:0] lut_962_select = {
                             in_data[66],
                             in_data[25],
                             in_data[741],
                             in_data[296],
                             in_data[239],
                             in_data[5]};
    
    wire lut_962_out = lut_962_table[lut_962_select];
    
    generate
    if ( USE_REG ) begin : ff_962
        reg   lut_962_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_962_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_962_ff <= lut_962_out;
            end
        end
        
        assign out_data[962] = lut_962_ff;
    end
    else begin : no_ff_962
        assign out_data[962] = lut_962_out;
    end
    endgenerate
    
    
    
    // LUT : 963
    wire [63:0] lut_963_table = 64'b1111000011110000111111111111111110100000100000001111111111111111;
    wire [5:0] lut_963_select = {
                             in_data[148],
                             in_data[412],
                             in_data[781],
                             in_data[525],
                             in_data[32],
                             in_data[307]};
    
    wire lut_963_out = lut_963_table[lut_963_select];
    
    generate
    if ( USE_REG ) begin : ff_963
        reg   lut_963_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_963_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_963_ff <= lut_963_out;
            end
        end
        
        assign out_data[963] = lut_963_ff;
    end
    else begin : no_ff_963
        assign out_data[963] = lut_963_out;
    end
    endgenerate
    
    
    
    // LUT : 964
    wire [63:0] lut_964_table = 64'b1111111111101110111111111110111100110000111000000011000011100000;
    wire [5:0] lut_964_select = {
                             in_data[184],
                             in_data[532],
                             in_data[514],
                             in_data[72],
                             in_data[329],
                             in_data[612]};
    
    wire lut_964_out = lut_964_table[lut_964_select];
    
    generate
    if ( USE_REG ) begin : ff_964
        reg   lut_964_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_964_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_964_ff <= lut_964_out;
            end
        end
        
        assign out_data[964] = lut_964_ff;
    end
    else begin : no_ff_964
        assign out_data[964] = lut_964_out;
    end
    endgenerate
    
    
    
    // LUT : 965
    wire [63:0] lut_965_table = 64'b0000010100010101000000000000000000000101000001010000000000000001;
    wire [5:0] lut_965_select = {
                             in_data[343],
                             in_data[607],
                             in_data[107],
                             in_data[176],
                             in_data[619],
                             in_data[146]};
    
    wire lut_965_out = lut_965_table[lut_965_select];
    
    generate
    if ( USE_REG ) begin : ff_965
        reg   lut_965_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_965_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_965_ff <= lut_965_out;
            end
        end
        
        assign out_data[965] = lut_965_ff;
    end
    else begin : no_ff_965
        assign out_data[965] = lut_965_out;
    end
    endgenerate
    
    
    
    // LUT : 966
    wire [63:0] lut_966_table = 64'b0111111101111111000000000011001100000000000000000000000000110011;
    wire [5:0] lut_966_select = {
                             in_data[435],
                             in_data[625],
                             in_data[485],
                             in_data[645],
                             in_data[469],
                             in_data[194]};
    
    wire lut_966_out = lut_966_table[lut_966_select];
    
    generate
    if ( USE_REG ) begin : ff_966
        reg   lut_966_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_966_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_966_ff <= lut_966_out;
            end
        end
        
        assign out_data[966] = lut_966_ff;
    end
    else begin : no_ff_966
        assign out_data[966] = lut_966_out;
    end
    endgenerate
    
    
    
    // LUT : 967
    wire [63:0] lut_967_table = 64'b0101011101010101010101110101010101000100010001000101010001010100;
    wire [5:0] lut_967_select = {
                             in_data[556],
                             in_data[472],
                             in_data[584],
                             in_data[319],
                             in_data[261],
                             in_data[96]};
    
    wire lut_967_out = lut_967_table[lut_967_select];
    
    generate
    if ( USE_REG ) begin : ff_967
        reg   lut_967_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_967_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_967_ff <= lut_967_out;
            end
        end
        
        assign out_data[967] = lut_967_ff;
    end
    else begin : no_ff_967
        assign out_data[967] = lut_967_out;
    end
    endgenerate
    
    
    
    // LUT : 968
    wire [63:0] lut_968_table = 64'b1111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_968_select = {
                             in_data[589],
                             in_data[783],
                             in_data[166],
                             in_data[187],
                             in_data[424],
                             in_data[731]};
    
    wire lut_968_out = lut_968_table[lut_968_select];
    
    generate
    if ( USE_REG ) begin : ff_968
        reg   lut_968_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_968_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_968_ff <= lut_968_out;
            end
        end
        
        assign out_data[968] = lut_968_ff;
    end
    else begin : no_ff_968
        assign out_data[968] = lut_968_out;
    end
    endgenerate
    
    
    
    // LUT : 969
    wire [63:0] lut_969_table = 64'b0001111100001010010111110000101001011111000010100101111100001110;
    wire [5:0] lut_969_select = {
                             in_data[776],
                             in_data[647],
                             in_data[570],
                             in_data[407],
                             in_data[467],
                             in_data[547]};
    
    wire lut_969_out = lut_969_table[lut_969_select];
    
    generate
    if ( USE_REG ) begin : ff_969
        reg   lut_969_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_969_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_969_ff <= lut_969_out;
            end
        end
        
        assign out_data[969] = lut_969_ff;
    end
    else begin : no_ff_969
        assign out_data[969] = lut_969_out;
    end
    endgenerate
    
    
    
    // LUT : 970
    wire [63:0] lut_970_table = 64'b0000000000000000101010101111111100000000000000000000000011111111;
    wire [5:0] lut_970_select = {
                             in_data[233],
                             in_data[132],
                             in_data[174],
                             in_data[0],
                             in_data[4],
                             in_data[219]};
    
    wire lut_970_out = lut_970_table[lut_970_select];
    
    generate
    if ( USE_REG ) begin : ff_970
        reg   lut_970_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_970_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_970_ff <= lut_970_out;
            end
        end
        
        assign out_data[970] = lut_970_ff;
    end
    else begin : no_ff_970
        assign out_data[970] = lut_970_out;
    end
    endgenerate
    
    
    
    // LUT : 971
    wire [63:0] lut_971_table = 64'b1111000011001000111100101110100011110011111010101111001111101010;
    wire [5:0] lut_971_select = {
                             in_data[431],
                             in_data[48],
                             in_data[440],
                             in_data[269],
                             in_data[382],
                             in_data[211]};
    
    wire lut_971_out = lut_971_table[lut_971_select];
    
    generate
    if ( USE_REG ) begin : ff_971
        reg   lut_971_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_971_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_971_ff <= lut_971_out;
            end
        end
        
        assign out_data[971] = lut_971_ff;
    end
    else begin : no_ff_971
        assign out_data[971] = lut_971_out;
    end
    endgenerate
    
    
    
    // LUT : 972
    wire [63:0] lut_972_table = 64'b1111111111111111111111111110111011111111111111111100110011001100;
    wire [5:0] lut_972_select = {
                             in_data[738],
                             in_data[710],
                             in_data[371],
                             in_data[20],
                             in_data[315],
                             in_data[213]};
    
    wire lut_972_out = lut_972_table[lut_972_select];
    
    generate
    if ( USE_REG ) begin : ff_972
        reg   lut_972_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_972_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_972_ff <= lut_972_out;
            end
        end
        
        assign out_data[972] = lut_972_ff;
    end
    else begin : no_ff_972
        assign out_data[972] = lut_972_out;
    end
    endgenerate
    
    
    
    // LUT : 973
    wire [63:0] lut_973_table = 64'b1111111111111111101010101110101011111111111111111010101010101010;
    wire [5:0] lut_973_select = {
                             in_data[644],
                             in_data[317],
                             in_data[295],
                             in_data[698],
                             in_data[53],
                             in_data[286]};
    
    wire lut_973_out = lut_973_table[lut_973_select];
    
    generate
    if ( USE_REG ) begin : ff_973
        reg   lut_973_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_973_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_973_ff <= lut_973_out;
            end
        end
        
        assign out_data[973] = lut_973_ff;
    end
    else begin : no_ff_973
        assign out_data[973] = lut_973_out;
    end
    endgenerate
    
    
    
    // LUT : 974
    wire [63:0] lut_974_table = 64'b0000000011111111000000000011011100000000111111110000000011001100;
    wire [5:0] lut_974_select = {
                             in_data[409],
                             in_data[419],
                             in_data[459],
                             in_data[669],
                             in_data[684],
                             in_data[585]};
    
    wire lut_974_out = lut_974_table[lut_974_select];
    
    generate
    if ( USE_REG ) begin : ff_974
        reg   lut_974_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_974_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_974_ff <= lut_974_out;
            end
        end
        
        assign out_data[974] = lut_974_ff;
    end
    else begin : no_ff_974
        assign out_data[974] = lut_974_out;
    end
    endgenerate
    
    
    
    // LUT : 975
    wire [63:0] lut_975_table = 64'b1111111100000000111111110000000011111111000000011111111100000000;
    wire [5:0] lut_975_select = {
                             in_data[775],
                             in_data[365],
                             in_data[359],
                             in_data[670],
                             in_data[423],
                             in_data[202]};
    
    wire lut_975_out = lut_975_table[lut_975_select];
    
    generate
    if ( USE_REG ) begin : ff_975
        reg   lut_975_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_975_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_975_ff <= lut_975_out;
            end
        end
        
        assign out_data[975] = lut_975_ff;
    end
    else begin : no_ff_975
        assign out_data[975] = lut_975_out;
    end
    endgenerate
    
    
    
    // LUT : 976
    wire [63:0] lut_976_table = 64'b1111111111111111110111011111111111111111111111110000000010001000;
    wire [5:0] lut_976_select = {
                             in_data[287],
                             in_data[341],
                             in_data[249],
                             in_data[112],
                             in_data[601],
                             in_data[388]};
    
    wire lut_976_out = lut_976_table[lut_976_select];
    
    generate
    if ( USE_REG ) begin : ff_976
        reg   lut_976_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_976_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_976_ff <= lut_976_out;
            end
        end
        
        assign out_data[976] = lut_976_ff;
    end
    else begin : no_ff_976
        assign out_data[976] = lut_976_out;
    end
    endgenerate
    
    
    
    // LUT : 977
    wire [63:0] lut_977_table = 64'b0000000001010101000000000101010000000000111111110000000011111111;
    wire [5:0] lut_977_select = {
                             in_data[492],
                             in_data[503],
                             in_data[411],
                             in_data[450],
                             in_data[34],
                             in_data[665]};
    
    wire lut_977_out = lut_977_table[lut_977_select];
    
    generate
    if ( USE_REG ) begin : ff_977
        reg   lut_977_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_977_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_977_ff <= lut_977_out;
            end
        end
        
        assign out_data[977] = lut_977_ff;
    end
    else begin : no_ff_977
        assign out_data[977] = lut_977_out;
    end
    endgenerate
    
    
    
    // LUT : 978
    wire [63:0] lut_978_table = 64'b1111111100000100111111110000010011111101010001011111110101000101;
    wire [5:0] lut_978_select = {
                             in_data[268],
                             in_data[560],
                             in_data[313],
                             in_data[175],
                             in_data[661],
                             in_data[283]};
    
    wire lut_978_out = lut_978_table[lut_978_select];
    
    generate
    if ( USE_REG ) begin : ff_978
        reg   lut_978_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_978_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_978_ff <= lut_978_out;
            end
        end
        
        assign out_data[978] = lut_978_ff;
    end
    else begin : no_ff_978
        assign out_data[978] = lut_978_out;
    end
    endgenerate
    
    
    
    // LUT : 979
    wire [63:0] lut_979_table = 64'b1111111111111111111111111111111011111111111000001111100011000000;
    wire [5:0] lut_979_select = {
                             in_data[515],
                             in_data[636],
                             in_data[385],
                             in_data[578],
                             in_data[756],
                             in_data[91]};
    
    wire lut_979_out = lut_979_table[lut_979_select];
    
    generate
    if ( USE_REG ) begin : ff_979
        reg   lut_979_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_979_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_979_ff <= lut_979_out;
            end
        end
        
        assign out_data[979] = lut_979_ff;
    end
    else begin : no_ff_979
        assign out_data[979] = lut_979_out;
    end
    endgenerate
    
    
    
    // LUT : 980
    wire [63:0] lut_980_table = 64'b1110100010000000111010001000000011111111111110111111111111111011;
    wire [5:0] lut_980_select = {
                             in_data[403],
                             in_data[506],
                             in_data[217],
                             in_data[133],
                             in_data[162],
                             in_data[263]};
    
    wire lut_980_out = lut_980_table[lut_980_select];
    
    generate
    if ( USE_REG ) begin : ff_980
        reg   lut_980_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_980_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_980_ff <= lut_980_out;
            end
        end
        
        assign out_data[980] = lut_980_ff;
    end
    else begin : no_ff_980
        assign out_data[980] = lut_980_out;
    end
    endgenerate
    
    
    
    // LUT : 981
    wire [63:0] lut_981_table = 64'b1111111111111111111111111111111111111111111111111111111100000000;
    wire [5:0] lut_981_select = {
                             in_data[487],
                             in_data[445],
                             in_data[157],
                             in_data[332],
                             in_data[753],
                             in_data[422]};
    
    wire lut_981_out = lut_981_table[lut_981_select];
    
    generate
    if ( USE_REG ) begin : ff_981
        reg   lut_981_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_981_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_981_ff <= lut_981_out;
            end
        end
        
        assign out_data[981] = lut_981_ff;
    end
    else begin : no_ff_981
        assign out_data[981] = lut_981_out;
    end
    endgenerate
    
    
    
    // LUT : 982
    wire [63:0] lut_982_table = 64'b0000111100001111000011110000111100000000000011110000000000001111;
    wire [5:0] lut_982_select = {
                             in_data[766],
                             in_data[46],
                             in_data[439],
                             in_data[415],
                             in_data[505],
                             in_data[30]};
    
    wire lut_982_out = lut_982_table[lut_982_select];
    
    generate
    if ( USE_REG ) begin : ff_982
        reg   lut_982_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_982_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_982_ff <= lut_982_out;
            end
        end
        
        assign out_data[982] = lut_982_ff;
    end
    else begin : no_ff_982
        assign out_data[982] = lut_982_out;
    end
    endgenerate
    
    
    
    // LUT : 983
    wire [63:0] lut_983_table = 64'b1111111111111111111111111111111111111111111111111110111011101110;
    wire [5:0] lut_983_select = {
                             in_data[565],
                             in_data[720],
                             in_data[526],
                             in_data[138],
                             in_data[554],
                             in_data[721]};
    
    wire lut_983_out = lut_983_table[lut_983_select];
    
    generate
    if ( USE_REG ) begin : ff_983
        reg   lut_983_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_983_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_983_ff <= lut_983_out;
            end
        end
        
        assign out_data[983] = lut_983_ff;
    end
    else begin : no_ff_983
        assign out_data[983] = lut_983_out;
    end
    endgenerate
    
    
    
    // LUT : 984
    wire [63:0] lut_984_table = 64'b1111111111101110111111111110111111101111111011101110111111101110;
    wire [5:0] lut_984_select = {
                             in_data[479],
                             in_data[35],
                             in_data[676],
                             in_data[311],
                             in_data[651],
                             in_data[404]};
    
    wire lut_984_out = lut_984_table[lut_984_select];
    
    generate
    if ( USE_REG ) begin : ff_984
        reg   lut_984_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_984_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_984_ff <= lut_984_out;
            end
        end
        
        assign out_data[984] = lut_984_ff;
    end
    else begin : no_ff_984
        assign out_data[984] = lut_984_out;
    end
    endgenerate
    
    
    
    // LUT : 985
    wire [63:0] lut_985_table = 64'b0000000000000000000000000000000000111011001110110000001000000010;
    wire [5:0] lut_985_select = {
                             in_data[723],
                             in_data[442],
                             in_data[2],
                             in_data[192],
                             in_data[255],
                             in_data[99]};
    
    wire lut_985_out = lut_985_table[lut_985_select];
    
    generate
    if ( USE_REG ) begin : ff_985
        reg   lut_985_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_985_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_985_ff <= lut_985_out;
            end
        end
        
        assign out_data[985] = lut_985_ff;
    end
    else begin : no_ff_985
        assign out_data[985] = lut_985_out;
    end
    endgenerate
    
    
    
    // LUT : 986
    wire [63:0] lut_986_table = 64'b1111111111111111110011001100110011111111111111111100110011001100;
    wire [5:0] lut_986_select = {
                             in_data[655],
                             in_data[123],
                             in_data[83],
                             in_data[690],
                             in_data[591],
                             in_data[726]};
    
    wire lut_986_out = lut_986_table[lut_986_select];
    
    generate
    if ( USE_REG ) begin : ff_986
        reg   lut_986_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_986_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_986_ff <= lut_986_out;
            end
        end
        
        assign out_data[986] = lut_986_ff;
    end
    else begin : no_ff_986
        assign out_data[986] = lut_986_out;
    end
    endgenerate
    
    
    
    // LUT : 987
    wire [63:0] lut_987_table = 64'b1110111011101110111111101111111110101010100011001000100010001000;
    wire [5:0] lut_987_select = {
                             in_data[353],
                             in_data[267],
                             in_data[364],
                             in_data[476],
                             in_data[209],
                             in_data[717]};
    
    wire lut_987_out = lut_987_table[lut_987_select];
    
    generate
    if ( USE_REG ) begin : ff_987
        reg   lut_987_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_987_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_987_ff <= lut_987_out;
            end
        end
        
        assign out_data[987] = lut_987_ff;
    end
    else begin : no_ff_987
        assign out_data[987] = lut_987_out;
    end
    endgenerate
    
    
    
    // LUT : 988
    wire [63:0] lut_988_table = 64'b1111001111110000111100111111001011110011111100101111001011110010;
    wire [5:0] lut_988_select = {
                             in_data[534],
                             in_data[393],
                             in_data[673],
                             in_data[681],
                             in_data[23],
                             in_data[51]};
    
    wire lut_988_out = lut_988_table[lut_988_select];
    
    generate
    if ( USE_REG ) begin : ff_988
        reg   lut_988_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_988_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_988_ff <= lut_988_out;
            end
        end
        
        assign out_data[988] = lut_988_ff;
    end
    else begin : no_ff_988
        assign out_data[988] = lut_988_out;
    end
    endgenerate
    
    
    
    // LUT : 989
    wire [63:0] lut_989_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_989_select = {
                             in_data[274],
                             in_data[74],
                             in_data[310],
                             in_data[615],
                             in_data[705],
                             in_data[410]};
    
    wire lut_989_out = lut_989_table[lut_989_select];
    
    generate
    if ( USE_REG ) begin : ff_989
        reg   lut_989_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_989_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_989_ff <= lut_989_out;
            end
        end
        
        assign out_data[989] = lut_989_ff;
    end
    else begin : no_ff_989
        assign out_data[989] = lut_989_out;
    end
    endgenerate
    
    
    
    // LUT : 990
    wire [63:0] lut_990_table = 64'b0000000000001111000000000000111111110000110111001111000011011100;
    wire [5:0] lut_990_select = {
                             in_data[594],
                             in_data[36],
                             in_data[320],
                             in_data[294],
                             in_data[545],
                             in_data[251]};
    
    wire lut_990_out = lut_990_table[lut_990_select];
    
    generate
    if ( USE_REG ) begin : ff_990
        reg   lut_990_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_990_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_990_ff <= lut_990_out;
            end
        end
        
        assign out_data[990] = lut_990_ff;
    end
    else begin : no_ff_990
        assign out_data[990] = lut_990_out;
    end
    endgenerate
    
    
    
    // LUT : 991
    wire [63:0] lut_991_table = 64'b1100110101001100111011111110111111001101010011001110111111101111;
    wire [5:0] lut_991_select = {
                             in_data[109],
                             in_data[379],
                             in_data[417],
                             in_data[163],
                             in_data[713],
                             in_data[273]};
    
    wire lut_991_out = lut_991_table[lut_991_select];
    
    generate
    if ( USE_REG ) begin : ff_991
        reg   lut_991_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_991_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_991_ff <= lut_991_out;
            end
        end
        
        assign out_data[991] = lut_991_ff;
    end
    else begin : no_ff_991
        assign out_data[991] = lut_991_out;
    end
    endgenerate
    
    
    
    // LUT : 992
    wire [63:0] lut_992_table = 64'b0001000100000000000100010000000011111111010001001111111101000000;
    wire [5:0] lut_992_select = {
                             in_data[256],
                             in_data[169],
                             in_data[321],
                             in_data[140],
                             in_data[355],
                             in_data[230]};
    
    wire lut_992_out = lut_992_table[lut_992_select];
    
    generate
    if ( USE_REG ) begin : ff_992
        reg   lut_992_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_992_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_992_ff <= lut_992_out;
            end
        end
        
        assign out_data[992] = lut_992_ff;
    end
    else begin : no_ff_992
        assign out_data[992] = lut_992_out;
    end
    endgenerate
    
    
    
    // LUT : 993
    wire [63:0] lut_993_table = 64'b1111111100110011111111110011001111111111000000100111111100000010;
    wire [5:0] lut_993_select = {
                             in_data[562],
                             in_data[701],
                             in_data[386],
                             in_data[727],
                             in_data[555],
                             in_data[730]};
    
    wire lut_993_out = lut_993_table[lut_993_select];
    
    generate
    if ( USE_REG ) begin : ff_993
        reg   lut_993_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_993_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_993_ff <= lut_993_out;
            end
        end
        
        assign out_data[993] = lut_993_ff;
    end
    else begin : no_ff_993
        assign out_data[993] = lut_993_out;
    end
    endgenerate
    
    
    
    // LUT : 994
    wire [63:0] lut_994_table = 64'b1111111111111111010101010000000011111111111111110101010100000000;
    wire [5:0] lut_994_select = {
                             in_data[779],
                             in_data[190],
                             in_data[304],
                             in_data[116],
                             in_data[448],
                             in_data[610]};
    
    wire lut_994_out = lut_994_table[lut_994_select];
    
    generate
    if ( USE_REG ) begin : ff_994
        reg   lut_994_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_994_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_994_ff <= lut_994_out;
            end
        end
        
        assign out_data[994] = lut_994_ff;
    end
    else begin : no_ff_994
        assign out_data[994] = lut_994_out;
    end
    endgenerate
    
    
    
    // LUT : 995
    wire [63:0] lut_995_table = 64'b0000111100000010111111110000111110001111000011101110111100001111;
    wire [5:0] lut_995_select = {
                             in_data[142],
                             in_data[481],
                             in_data[368],
                             in_data[463],
                             in_data[58],
                             in_data[497]};
    
    wire lut_995_out = lut_995_table[lut_995_select];
    
    generate
    if ( USE_REG ) begin : ff_995
        reg   lut_995_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_995_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_995_ff <= lut_995_out;
            end
        end
        
        assign out_data[995] = lut_995_ff;
    end
    else begin : no_ff_995
        assign out_data[995] = lut_995_out;
    end
    endgenerate
    
    
    
    // LUT : 996
    wire [63:0] lut_996_table = 64'b0000000011111111000000001111111100000000110111010000000011111111;
    wire [5:0] lut_996_select = {
                             in_data[675],
                             in_data[61],
                             in_data[453],
                             in_data[19],
                             in_data[643],
                             in_data[752]};
    
    wire lut_996_out = lut_996_table[lut_996_select];
    
    generate
    if ( USE_REG ) begin : ff_996
        reg   lut_996_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_996_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_996_ff <= lut_996_out;
            end
        end
        
        assign out_data[996] = lut_996_ff;
    end
    else begin : no_ff_996
        assign out_data[996] = lut_996_out;
    end
    endgenerate
    
    
    
    // LUT : 997
    wire [63:0] lut_997_table = 64'b0000000000000100110000001111000011110100111111011111000011111100;
    wire [5:0] lut_997_select = {
                             in_data[563],
                             in_data[272],
                             in_data[557],
                             in_data[301],
                             in_data[627],
                             in_data[735]};
    
    wire lut_997_out = lut_997_table[lut_997_select];
    
    generate
    if ( USE_REG ) begin : ff_997
        reg   lut_997_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_997_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_997_ff <= lut_997_out;
            end
        end
        
        assign out_data[997] = lut_997_ff;
    end
    else begin : no_ff_997
        assign out_data[997] = lut_997_out;
    end
    endgenerate
    
    
    
    // LUT : 998
    wire [63:0] lut_998_table = 64'b0011001111111111001100111111011100110011111111110011001100110011;
    wire [5:0] lut_998_select = {
                             in_data[220],
                             in_data[156],
                             in_data[344],
                             in_data[200],
                             in_data[186],
                             in_data[765]};
    
    wire lut_998_out = lut_998_table[lut_998_select];
    
    generate
    if ( USE_REG ) begin : ff_998
        reg   lut_998_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_998_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_998_ff <= lut_998_out;
            end
        end
        
        assign out_data[998] = lut_998_ff;
    end
    else begin : no_ff_998
        assign out_data[998] = lut_998_out;
    end
    endgenerate
    
    
    
    // LUT : 999
    wire [63:0] lut_999_table = 64'b1111110011111100110000001100000011111100111111001100000011000000;
    wire [5:0] lut_999_select = {
                             in_data[559],
                             in_data[443],
                             in_data[227],
                             in_data[572],
                             in_data[548],
                             in_data[590]};
    
    wire lut_999_out = lut_999_table[lut_999_select];
    
    generate
    if ( USE_REG ) begin : ff_999
        reg   lut_999_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_999_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_999_ff <= lut_999_out;
            end
        end
        
        assign out_data[999] = lut_999_ff;
    end
    else begin : no_ff_999
        assign out_data[999] = lut_999_out;
    end
    endgenerate
    
    
    
    // LUT : 1000
    wire [63:0] lut_1000_table = 64'b1111001101110000001000101010001011110011111100011010101010101010;
    wire [5:0] lut_1000_select = {
                             in_data[37],
                             in_data[523],
                             in_data[188],
                             in_data[518],
                             in_data[305],
                             in_data[580]};
    
    wire lut_1000_out = lut_1000_table[lut_1000_select];
    
    generate
    if ( USE_REG ) begin : ff_1000
        reg   lut_1000_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1000_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1000_ff <= lut_1000_out;
            end
        end
        
        assign out_data[1000] = lut_1000_ff;
    end
    else begin : no_ff_1000
        assign out_data[1000] = lut_1000_out;
    end
    endgenerate
    
    
    
    // LUT : 1001
    wire [63:0] lut_1001_table = 64'b0001001100110011001000100011001100000011001100110010001000110011;
    wire [5:0] lut_1001_select = {
                             in_data[749],
                             in_data[264],
                             in_data[474],
                             in_data[401],
                             in_data[324],
                             in_data[318]};
    
    wire lut_1001_out = lut_1001_table[lut_1001_select];
    
    generate
    if ( USE_REG ) begin : ff_1001
        reg   lut_1001_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1001_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1001_ff <= lut_1001_out;
            end
        end
        
        assign out_data[1001] = lut_1001_ff;
    end
    else begin : no_ff_1001
        assign out_data[1001] = lut_1001_out;
    end
    endgenerate
    
    
    
    // LUT : 1002
    wire [63:0] lut_1002_table = 64'b1000111110101111101011111010111111111010101110101111101010111010;
    wire [5:0] lut_1002_select = {
                             in_data[438],
                             in_data[671],
                             in_data[361],
                             in_data[495],
                             in_data[432],
                             in_data[266]};
    
    wire lut_1002_out = lut_1002_table[lut_1002_select];
    
    generate
    if ( USE_REG ) begin : ff_1002
        reg   lut_1002_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1002_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1002_ff <= lut_1002_out;
            end
        end
        
        assign out_data[1002] = lut_1002_ff;
    end
    else begin : no_ff_1002
        assign out_data[1002] = lut_1002_out;
    end
    endgenerate
    
    
    
    // LUT : 1003
    wire [63:0] lut_1003_table = 64'b0000000010111111111111110010001100001000101011111100110000000011;
    wire [5:0] lut_1003_select = {
                             in_data[648],
                             in_data[402],
                             in_data[662],
                             in_data[656],
                             in_data[325],
                             in_data[672]};
    
    wire lut_1003_out = lut_1003_table[lut_1003_select];
    
    generate
    if ( USE_REG ) begin : ff_1003
        reg   lut_1003_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1003_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1003_ff <= lut_1003_out;
            end
        end
        
        assign out_data[1003] = lut_1003_ff;
    end
    else begin : no_ff_1003
        assign out_data[1003] = lut_1003_out;
    end
    endgenerate
    
    
    
    // LUT : 1004
    wire [63:0] lut_1004_table = 64'b0000000000000011000000000000001101110011111100111111011111110011;
    wire [5:0] lut_1004_select = {
                             in_data[430],
                             in_data[338],
                             in_data[456],
                             in_data[659],
                             in_data[541],
                             in_data[136]};
    
    wire lut_1004_out = lut_1004_table[lut_1004_select];
    
    generate
    if ( USE_REG ) begin : ff_1004
        reg   lut_1004_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1004_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1004_ff <= lut_1004_out;
            end
        end
        
        assign out_data[1004] = lut_1004_ff;
    end
    else begin : no_ff_1004
        assign out_data[1004] = lut_1004_out;
    end
    endgenerate
    
    
    
    // LUT : 1005
    wire [63:0] lut_1005_table = 64'b1110101011101010111110111111101011101010111010101111101111101010;
    wire [5:0] lut_1005_select = {
                             in_data[144],
                             in_data[300],
                             in_data[285],
                             in_data[494],
                             in_data[356],
                             in_data[553]};
    
    wire lut_1005_out = lut_1005_table[lut_1005_select];
    
    generate
    if ( USE_REG ) begin : ff_1005
        reg   lut_1005_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1005_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1005_ff <= lut_1005_out;
            end
        end
        
        assign out_data[1005] = lut_1005_ff;
    end
    else begin : no_ff_1005
        assign out_data[1005] = lut_1005_out;
    end
    endgenerate
    
    
    
    // LUT : 1006
    wire [63:0] lut_1006_table = 64'b1111010011110101111101011111010111110000111101011111000111110101;
    wire [5:0] lut_1006_select = {
                             in_data[778],
                             in_data[508],
                             in_data[704],
                             in_data[745],
                             in_data[12],
                             in_data[270]};
    
    wire lut_1006_out = lut_1006_table[lut_1006_select];
    
    generate
    if ( USE_REG ) begin : ff_1006
        reg   lut_1006_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1006_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1006_ff <= lut_1006_out;
            end
        end
        
        assign out_data[1006] = lut_1006_ff;
    end
    else begin : no_ff_1006
        assign out_data[1006] = lut_1006_out;
    end
    endgenerate
    
    
    
    // LUT : 1007
    wire [63:0] lut_1007_table = 64'b0000000000000000000000000000000011111111111110001111111111101111;
    wire [5:0] lut_1007_select = {
                             in_data[689],
                             in_data[739],
                             in_data[677],
                             in_data[236],
                             in_data[15],
                             in_data[52]};
    
    wire lut_1007_out = lut_1007_table[lut_1007_select];
    
    generate
    if ( USE_REG ) begin : ff_1007
        reg   lut_1007_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1007_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1007_ff <= lut_1007_out;
            end
        end
        
        assign out_data[1007] = lut_1007_ff;
    end
    else begin : no_ff_1007
        assign out_data[1007] = lut_1007_out;
    end
    endgenerate
    
    
    
    // LUT : 1008
    wire [63:0] lut_1008_table = 64'b1100110010001100110011001000110011001100000011001100110010001100;
    wire [5:0] lut_1008_select = {
                             in_data[31],
                             in_data[641],
                             in_data[105],
                             in_data[247],
                             in_data[381],
                             in_data[782]};
    
    wire lut_1008_out = lut_1008_table[lut_1008_select];
    
    generate
    if ( USE_REG ) begin : ff_1008
        reg   lut_1008_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1008_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1008_ff <= lut_1008_out;
            end
        end
        
        assign out_data[1008] = lut_1008_ff;
    end
    else begin : no_ff_1008
        assign out_data[1008] = lut_1008_out;
    end
    endgenerate
    
    
    
    // LUT : 1009
    wire [63:0] lut_1009_table = 64'b0111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_1009_select = {
                             in_data[245],
                             in_data[466],
                             in_data[632],
                             in_data[158],
                             in_data[168],
                             in_data[151]};
    
    wire lut_1009_out = lut_1009_table[lut_1009_select];
    
    generate
    if ( USE_REG ) begin : ff_1009
        reg   lut_1009_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1009_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1009_ff <= lut_1009_out;
            end
        end
        
        assign out_data[1009] = lut_1009_ff;
    end
    else begin : no_ff_1009
        assign out_data[1009] = lut_1009_out;
    end
    endgenerate
    
    
    
    // LUT : 1010
    wire [63:0] lut_1010_table = 64'b1111111111111111111111111111111111110000111100001111000011110000;
    wire [5:0] lut_1010_select = {
                             in_data[653],
                             in_data[759],
                             in_data[281],
                             in_data[288],
                             in_data[6],
                             in_data[85]};
    
    wire lut_1010_out = lut_1010_table[lut_1010_select];
    
    generate
    if ( USE_REG ) begin : ff_1010
        reg   lut_1010_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1010_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1010_ff <= lut_1010_out;
            end
        end
        
        assign out_data[1010] = lut_1010_ff;
    end
    else begin : no_ff_1010
        assign out_data[1010] = lut_1010_out;
    end
    endgenerate
    
    
    
    // LUT : 1011
    wire [63:0] lut_1011_table = 64'b1111111111111111110011001101110111111111111111110000000000000000;
    wire [5:0] lut_1011_select = {
                             in_data[748],
                             in_data[183],
                             in_data[291],
                             in_data[10],
                             in_data[524],
                             in_data[384]};
    
    wire lut_1011_out = lut_1011_table[lut_1011_select];
    
    generate
    if ( USE_REG ) begin : ff_1011
        reg   lut_1011_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1011_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1011_ff <= lut_1011_out;
            end
        end
        
        assign out_data[1011] = lut_1011_ff;
    end
    else begin : no_ff_1011
        assign out_data[1011] = lut_1011_out;
    end
    endgenerate
    
    
    
    // LUT : 1012
    wire [63:0] lut_1012_table = 64'b0000000000000001000000000011001100000000000000000000000000010011;
    wire [5:0] lut_1012_select = {
                             in_data[57],
                             in_data[529],
                             in_data[124],
                             in_data[29],
                             in_data[510],
                             in_data[640]};
    
    wire lut_1012_out = lut_1012_table[lut_1012_select];
    
    generate
    if ( USE_REG ) begin : ff_1012
        reg   lut_1012_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1012_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1012_ff <= lut_1012_out;
            end
        end
        
        assign out_data[1012] = lut_1012_ff;
    end
    else begin : no_ff_1012
        assign out_data[1012] = lut_1012_out;
    end
    endgenerate
    
    
    
    // LUT : 1013
    wire [63:0] lut_1013_table = 64'b1000100010001100100010001000110011011101111111111101110111111111;
    wire [5:0] lut_1013_select = {
                             in_data[493],
                             in_data[108],
                             in_data[606],
                             in_data[279],
                             in_data[303],
                             in_data[351]};
    
    wire lut_1013_out = lut_1013_table[lut_1013_select];
    
    generate
    if ( USE_REG ) begin : ff_1013
        reg   lut_1013_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1013_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1013_ff <= lut_1013_out;
            end
        end
        
        assign out_data[1013] = lut_1013_ff;
    end
    else begin : no_ff_1013
        assign out_data[1013] = lut_1013_out;
    end
    endgenerate
    
    
    
    // LUT : 1014
    wire [63:0] lut_1014_table = 64'b1111101111111011011100110101001011110011111110110101001101010000;
    wire [5:0] lut_1014_select = {
                             in_data[362],
                             in_data[736],
                             in_data[638],
                             in_data[290],
                             in_data[688],
                             in_data[265]};
    
    wire lut_1014_out = lut_1014_table[lut_1014_select];
    
    generate
    if ( USE_REG ) begin : ff_1014
        reg   lut_1014_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1014_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1014_ff <= lut_1014_out;
            end
        end
        
        assign out_data[1014] = lut_1014_ff;
    end
    else begin : no_ff_1014
        assign out_data[1014] = lut_1014_out;
    end
    endgenerate
    
    
    
    // LUT : 1015
    wire [63:0] lut_1015_table = 64'b1100110011000000110000001100000011001100110011001111110011111100;
    wire [5:0] lut_1015_select = {
                             in_data[629],
                             in_data[605],
                             in_data[342],
                             in_data[289],
                             in_data[354],
                             in_data[13]};
    
    wire lut_1015_out = lut_1015_table[lut_1015_select];
    
    generate
    if ( USE_REG ) begin : ff_1015
        reg   lut_1015_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1015_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1015_ff <= lut_1015_out;
            end
        end
        
        assign out_data[1015] = lut_1015_ff;
    end
    else begin : no_ff_1015
        assign out_data[1015] = lut_1015_out;
    end
    endgenerate
    
    
    
    // LUT : 1016
    wire [63:0] lut_1016_table = 64'b0000000000000000000100000011001111001100000000001011001110110011;
    wire [5:0] lut_1016_select = {
                             in_data[185],
                             in_data[436],
                             in_data[623],
                             in_data[366],
                             in_data[491],
                             in_data[418]};
    
    wire lut_1016_out = lut_1016_table[lut_1016_select];
    
    generate
    if ( USE_REG ) begin : ff_1016
        reg   lut_1016_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1016_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1016_ff <= lut_1016_out;
            end
        end
        
        assign out_data[1016] = lut_1016_ff;
    end
    else begin : no_ff_1016
        assign out_data[1016] = lut_1016_out;
    end
    endgenerate
    
    
    
    // LUT : 1017
    wire [63:0] lut_1017_table = 64'b1100000001000000000000001100110011100000000000001110000011111100;
    wire [5:0] lut_1017_select = {
                             in_data[692],
                             in_data[539],
                             in_data[101],
                             in_data[240],
                             in_data[746],
                             in_data[308]};
    
    wire lut_1017_out = lut_1017_table[lut_1017_select];
    
    generate
    if ( USE_REG ) begin : ff_1017
        reg   lut_1017_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1017_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1017_ff <= lut_1017_out;
            end
        end
        
        assign out_data[1017] = lut_1017_ff;
    end
    else begin : no_ff_1017
        assign out_data[1017] = lut_1017_out;
    end
    endgenerate
    
    
    
    // LUT : 1018
    wire [63:0] lut_1018_table = 64'b1111111111111111111111111000100011111111111111111111111110001000;
    wire [5:0] lut_1018_select = {
                             in_data[250],
                             in_data[126],
                             in_data[441],
                             in_data[8],
                             in_data[568],
                             in_data[154]};
    
    wire lut_1018_out = lut_1018_table[lut_1018_select];
    
    generate
    if ( USE_REG ) begin : ff_1018
        reg   lut_1018_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1018_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1018_ff <= lut_1018_out;
            end
        end
        
        assign out_data[1018] = lut_1018_ff;
    end
    else begin : no_ff_1018
        assign out_data[1018] = lut_1018_out;
    end
    endgenerate
    
    
    
    // LUT : 1019
    wire [63:0] lut_1019_table = 64'b1010101110101011101010111010101100001010000010100000101000001010;
    wire [5:0] lut_1019_select = {
                             in_data[551],
                             in_data[44],
                             in_data[1],
                             in_data[98],
                             in_data[218],
                             in_data[298]};
    
    wire lut_1019_out = lut_1019_table[lut_1019_select];
    
    generate
    if ( USE_REG ) begin : ff_1019
        reg   lut_1019_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1019_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1019_ff <= lut_1019_out;
            end
        end
        
        assign out_data[1019] = lut_1019_ff;
    end
    else begin : no_ff_1019
        assign out_data[1019] = lut_1019_out;
    end
    endgenerate
    
    
    
    // LUT : 1020
    wire [63:0] lut_1020_table = 64'b0000000000000000000000000000000000000000000000000001000100010001;
    wire [5:0] lut_1020_select = {
                             in_data[161],
                             in_data[770],
                             in_data[392],
                             in_data[24],
                             in_data[306],
                             in_data[191]};
    
    wire lut_1020_out = lut_1020_table[lut_1020_select];
    
    generate
    if ( USE_REG ) begin : ff_1020
        reg   lut_1020_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1020_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1020_ff <= lut_1020_out;
            end
        end
        
        assign out_data[1020] = lut_1020_ff;
    end
    else begin : no_ff_1020
        assign out_data[1020] = lut_1020_out;
    end
    endgenerate
    
    
    
    // LUT : 1021
    wire [63:0] lut_1021_table = 64'b1101010011010100110101001101010011010101110111001101110111010100;
    wire [5:0] lut_1021_select = {
                             in_data[737],
                             in_data[760],
                             in_data[498],
                             in_data[248],
                             in_data[374],
                             in_data[549]};
    
    wire lut_1021_out = lut_1021_table[lut_1021_select];
    
    generate
    if ( USE_REG ) begin : ff_1021
        reg   lut_1021_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1021_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1021_ff <= lut_1021_out;
            end
        end
        
        assign out_data[1021] = lut_1021_ff;
    end
    else begin : no_ff_1021
        assign out_data[1021] = lut_1021_out;
    end
    endgenerate
    
    
    
    // LUT : 1022
    wire [63:0] lut_1022_table = 64'b1100110011001100000000000000000011001100110011001100110011001100;
    wire [5:0] lut_1022_select = {
                             in_data[94],
                             in_data[634],
                             in_data[695],
                             in_data[276],
                             in_data[519],
                             in_data[42]};
    
    wire lut_1022_out = lut_1022_table[lut_1022_select];
    
    generate
    if ( USE_REG ) begin : ff_1022
        reg   lut_1022_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1022_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1022_ff <= lut_1022_out;
            end
        end
        
        assign out_data[1022] = lut_1022_ff;
    end
    else begin : no_ff_1022
        assign out_data[1022] = lut_1022_out;
    end
    endgenerate
    
    
    
    // LUT : 1023
    wire [63:0] lut_1023_table = 64'b0000110000000000110011011100110001001100010000001100110111001100;
    wire [5:0] lut_1023_select = {
                             in_data[334],
                             in_data[257],
                             in_data[397],
                             in_data[358],
                             in_data[462],
                             in_data[774]};
    
    wire lut_1023_out = lut_1023_table[lut_1023_select];
    
    generate
    if ( USE_REG ) begin : ff_1023
        reg   lut_1023_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1023_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1023_ff <= lut_1023_out;
            end
        end
        
        assign out_data[1023] = lut_1023_ff;
    end
    else begin : no_ff_1023
        assign out_data[1023] = lut_1023_out;
    end
    endgenerate
    
    
    
    // LUT : 1024
    wire [63:0] lut_1024_table = 64'b1111111111111111111111111111111111111111001100111111111100010001;
    wire [5:0] lut_1024_select = {
                             in_data[149],
                             in_data[309],
                             in_data[633],
                             in_data[561],
                             in_data[243],
                             in_data[678]};
    
    wire lut_1024_out = lut_1024_table[lut_1024_select];
    
    generate
    if ( USE_REG ) begin : ff_1024
        reg   lut_1024_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1024_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1024_ff <= lut_1024_out;
            end
        end
        
        assign out_data[1024] = lut_1024_ff;
    end
    else begin : no_ff_1024
        assign out_data[1024] = lut_1024_out;
    end
    endgenerate
    
    
    
    // LUT : 1025
    wire [63:0] lut_1025_table = 64'b0000000000000000000000000000000011111111010101011111111101010101;
    wire [5:0] lut_1025_select = {
                             in_data[125],
                             in_data[56],
                             in_data[221],
                             in_data[449],
                             in_data[363],
                             in_data[552]};
    
    wire lut_1025_out = lut_1025_table[lut_1025_select];
    
    generate
    if ( USE_REG ) begin : ff_1025
        reg   lut_1025_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1025_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1025_ff <= lut_1025_out;
            end
        end
        
        assign out_data[1025] = lut_1025_ff;
    end
    else begin : no_ff_1025
        assign out_data[1025] = lut_1025_out;
    end
    endgenerate
    
    
    
    // LUT : 1026
    wire [63:0] lut_1026_table = 64'b1111010011110100111111111111111111100100111001001111010111110100;
    wire [5:0] lut_1026_select = {
                             in_data[134],
                             in_data[620],
                             in_data[41],
                             in_data[718],
                             in_data[314],
                             in_data[520]};
    
    wire lut_1026_out = lut_1026_table[lut_1026_select];
    
    generate
    if ( USE_REG ) begin : ff_1026
        reg   lut_1026_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1026_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1026_ff <= lut_1026_out;
            end
        end
        
        assign out_data[1026] = lut_1026_ff;
    end
    else begin : no_ff_1026
        assign out_data[1026] = lut_1026_out;
    end
    endgenerate
    
    
    
    // LUT : 1027
    wire [63:0] lut_1027_table = 64'b0000111100001111000000110000001100001111000011110000001100000011;
    wire [5:0] lut_1027_select = {
                             in_data[62],
                             in_data[328],
                             in_data[639],
                             in_data[537],
                             in_data[348],
                             in_data[252]};
    
    wire lut_1027_out = lut_1027_table[lut_1027_select];
    
    generate
    if ( USE_REG ) begin : ff_1027
        reg   lut_1027_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1027_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1027_ff <= lut_1027_out;
            end
        end
        
        assign out_data[1027] = lut_1027_ff;
    end
    else begin : no_ff_1027
        assign out_data[1027] = lut_1027_out;
    end
    endgenerate
    
    
    
    // LUT : 1028
    wire [63:0] lut_1028_table = 64'b0011000000110000011100000111000000110000011100000111000011110001;
    wire [5:0] lut_1028_select = {
                             in_data[504],
                             in_data[75],
                             in_data[768],
                             in_data[598],
                             in_data[575],
                             in_data[77]};
    
    wire lut_1028_out = lut_1028_table[lut_1028_select];
    
    generate
    if ( USE_REG ) begin : ff_1028
        reg   lut_1028_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1028_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1028_ff <= lut_1028_out;
            end
        end
        
        assign out_data[1028] = lut_1028_ff;
    end
    else begin : no_ff_1028
        assign out_data[1028] = lut_1028_out;
    end
    endgenerate
    
    
    
    // LUT : 1029
    wire [63:0] lut_1029_table = 64'b0011001100110011001100110011001100000000000000000000000000000000;
    wire [5:0] lut_1029_select = {
                             in_data[378],
                             in_data[587],
                             in_data[60],
                             in_data[253],
                             in_data[719],
                             in_data[203]};
    
    wire lut_1029_out = lut_1029_table[lut_1029_select];
    
    generate
    if ( USE_REG ) begin : ff_1029
        reg   lut_1029_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1029_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1029_ff <= lut_1029_out;
            end
        end
        
        assign out_data[1029] = lut_1029_ff;
    end
    else begin : no_ff_1029
        assign out_data[1029] = lut_1029_out;
    end
    endgenerate
    
    
    
    // LUT : 1030
    wire [63:0] lut_1030_table = 64'b0101010101010000010101010101000001010101111100000101010101110101;
    wire [5:0] lut_1030_select = {
                             in_data[135],
                             in_data[399],
                             in_data[201],
                             in_data[666],
                             in_data[333],
                             in_data[376]};
    
    wire lut_1030_out = lut_1030_table[lut_1030_select];
    
    generate
    if ( USE_REG ) begin : ff_1030
        reg   lut_1030_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1030_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1030_ff <= lut_1030_out;
            end
        end
        
        assign out_data[1030] = lut_1030_ff;
    end
    else begin : no_ff_1030
        assign out_data[1030] = lut_1030_out;
    end
    endgenerate
    
    
    
    // LUT : 1031
    wire [63:0] lut_1031_table = 64'b1111111111110011111111111111111110100000101000001011001010110010;
    wire [5:0] lut_1031_select = {
                             in_data[207],
                             in_data[535],
                             in_data[198],
                             in_data[327],
                             in_data[223],
                             in_data[235]};
    
    wire lut_1031_out = lut_1031_table[lut_1031_select];
    
    generate
    if ( USE_REG ) begin : ff_1031
        reg   lut_1031_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1031_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1031_ff <= lut_1031_out;
            end
        end
        
        assign out_data[1031] = lut_1031_ff;
    end
    else begin : no_ff_1031
        assign out_data[1031] = lut_1031_out;
    end
    endgenerate
    
    
    
    // LUT : 1032
    wire [63:0] lut_1032_table = 64'b1111010111110100110100000100000011111101111111111111010011111101;
    wire [5:0] lut_1032_select = {
                             in_data[455],
                             in_data[722],
                             in_data[444],
                             in_data[103],
                             in_data[763],
                             in_data[69]};
    
    wire lut_1032_out = lut_1032_table[lut_1032_select];
    
    generate
    if ( USE_REG ) begin : ff_1032
        reg   lut_1032_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1032_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1032_ff <= lut_1032_out;
            end
        end
        
        assign out_data[1032] = lut_1032_ff;
    end
    else begin : no_ff_1032
        assign out_data[1032] = lut_1032_out;
    end
    endgenerate
    
    
    
    // LUT : 1033
    wire [63:0] lut_1033_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1033_select = {
                             in_data[160],
                             in_data[408],
                             in_data[702],
                             in_data[579],
                             in_data[400],
                             in_data[751]};
    
    wire lut_1033_out = lut_1033_table[lut_1033_select];
    
    generate
    if ( USE_REG ) begin : ff_1033
        reg   lut_1033_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1033_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1033_ff <= lut_1033_out;
            end
        end
        
        assign out_data[1033] = lut_1033_ff;
    end
    else begin : no_ff_1033
        assign out_data[1033] = lut_1033_out;
    end
    endgenerate
    
    
    
    // LUT : 1034
    wire [63:0] lut_1034_table = 64'b0000000000000000000000000001000100000000000000000000000000010001;
    wire [5:0] lut_1034_select = {
                             in_data[232],
                             in_data[744],
                             in_data[164],
                             in_data[14],
                             in_data[100],
                             in_data[667]};
    
    wire lut_1034_out = lut_1034_table[lut_1034_select];
    
    generate
    if ( USE_REG ) begin : ff_1034
        reg   lut_1034_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1034_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1034_ff <= lut_1034_out;
            end
        end
        
        assign out_data[1034] = lut_1034_ff;
    end
    else begin : no_ff_1034
        assign out_data[1034] = lut_1034_out;
    end
    endgenerate
    
    
    
    // LUT : 1035
    wire [63:0] lut_1035_table = 64'b1111111100110011001100110000001011111111001100110011001100000000;
    wire [5:0] lut_1035_select = {
                             in_data[533],
                             in_data[528],
                             in_data[260],
                             in_data[139],
                             in_data[567],
                             in_data[111]};
    
    wire lut_1035_out = lut_1035_table[lut_1035_select];
    
    generate
    if ( USE_REG ) begin : ff_1035
        reg   lut_1035_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1035_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1035_ff <= lut_1035_out;
            end
        end
        
        assign out_data[1035] = lut_1035_ff;
    end
    else begin : no_ff_1035
        assign out_data[1035] = lut_1035_out;
    end
    endgenerate
    
    
    
    // LUT : 1036
    wire [63:0] lut_1036_table = 64'b0000000000000000000000000000000011111111000000001111111111111111;
    wire [5:0] lut_1036_select = {
                             in_data[742],
                             in_data[337],
                             in_data[254],
                             in_data[59],
                             in_data[196],
                             in_data[49]};
    
    wire lut_1036_out = lut_1036_table[lut_1036_select];
    
    generate
    if ( USE_REG ) begin : ff_1036
        reg   lut_1036_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1036_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1036_ff <= lut_1036_out;
            end
        end
        
        assign out_data[1036] = lut_1036_ff;
    end
    else begin : no_ff_1036
        assign out_data[1036] = lut_1036_out;
    end
    endgenerate
    
    
    
    // LUT : 1037
    wire [63:0] lut_1037_table = 64'b1101111100001111110111110000111001011111000011111111111100000000;
    wire [5:0] lut_1037_select = {
                             in_data[170],
                             in_data[204],
                             in_data[189],
                             in_data[454],
                             in_data[729],
                             in_data[687]};
    
    wire lut_1037_out = lut_1037_table[lut_1037_select];
    
    generate
    if ( USE_REG ) begin : ff_1037
        reg   lut_1037_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1037_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1037_ff <= lut_1037_out;
            end
        end
        
        assign out_data[1037] = lut_1037_ff;
    end
    else begin : no_ff_1037
        assign out_data[1037] = lut_1037_out;
    end
    endgenerate
    
    
    
    // LUT : 1038
    wire [63:0] lut_1038_table = 64'b0000000000000000000000000000000000110000011100010011000001110001;
    wire [5:0] lut_1038_select = {
                             in_data[210],
                             in_data[39],
                             in_data[500],
                             in_data[544],
                             in_data[593],
                             in_data[95]};
    
    wire lut_1038_out = lut_1038_table[lut_1038_select];
    
    generate
    if ( USE_REG ) begin : ff_1038
        reg   lut_1038_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1038_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1038_ff <= lut_1038_out;
            end
        end
        
        assign out_data[1038] = lut_1038_ff;
    end
    else begin : no_ff_1038
        assign out_data[1038] = lut_1038_out;
    end
    endgenerate
    
    
    
    // LUT : 1039
    wire [63:0] lut_1039_table = 64'b1111111110101111111111111111111111111111111111111111111100000000;
    wire [5:0] lut_1039_select = {
                             in_data[150],
                             in_data[482],
                             in_data[275],
                             in_data[115],
                             in_data[613],
                             in_data[699]};
    
    wire lut_1039_out = lut_1039_table[lut_1039_select];
    
    generate
    if ( USE_REG ) begin : ff_1039
        reg   lut_1039_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1039_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1039_ff <= lut_1039_out;
            end
        end
        
        assign out_data[1039] = lut_1039_ff;
    end
    else begin : no_ff_1039
        assign out_data[1039] = lut_1039_out;
    end
    endgenerate
    
    
    
    // LUT : 1040
    wire [63:0] lut_1040_table = 64'b1111111111111111110011001100110011111111111111111111111111111111;
    wire [5:0] lut_1040_select = {
                             in_data[543],
                             in_data[706],
                             in_data[780],
                             in_data[87],
                             in_data[428],
                             in_data[703]};
    
    wire lut_1040_out = lut_1040_table[lut_1040_select];
    
    generate
    if ( USE_REG ) begin : ff_1040
        reg   lut_1040_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1040_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1040_ff <= lut_1040_out;
            end
        end
        
        assign out_data[1040] = lut_1040_ff;
    end
    else begin : no_ff_1040
        assign out_data[1040] = lut_1040_out;
    end
    endgenerate
    
    
    
    // LUT : 1041
    wire [63:0] lut_1041_table = 64'b1111111100000000111111111111111111101110000000001111111111111111;
    wire [5:0] lut_1041_select = {
                             in_data[756],
                             in_data[345],
                             in_data[396],
                             in_data[363],
                             in_data[542],
                             in_data[1]};
    
    wire lut_1041_out = lut_1041_table[lut_1041_select];
    
    generate
    if ( USE_REG ) begin : ff_1041
        reg   lut_1041_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1041_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1041_ff <= lut_1041_out;
            end
        end
        
        assign out_data[1041] = lut_1041_ff;
    end
    else begin : no_ff_1041
        assign out_data[1041] = lut_1041_out;
    end
    endgenerate
    
    
    
    // LUT : 1042
    wire [63:0] lut_1042_table = 64'b0000000000000000000000000000000000000000000011110000000000001111;
    wire [5:0] lut_1042_select = {
                             in_data[213],
                             in_data[336],
                             in_data[711],
                             in_data[566],
                             in_data[590],
                             in_data[504]};
    
    wire lut_1042_out = lut_1042_table[lut_1042_select];
    
    generate
    if ( USE_REG ) begin : ff_1042
        reg   lut_1042_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1042_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1042_ff <= lut_1042_out;
            end
        end
        
        assign out_data[1042] = lut_1042_ff;
    end
    else begin : no_ff_1042
        assign out_data[1042] = lut_1042_out;
    end
    endgenerate
    
    
    
    // LUT : 1043
    wire [63:0] lut_1043_table = 64'b1111111111111111111111111111111101010101000100010100010000000000;
    wire [5:0] lut_1043_select = {
                             in_data[154],
                             in_data[669],
                             in_data[603],
                             in_data[89],
                             in_data[61],
                             in_data[326]};
    
    wire lut_1043_out = lut_1043_table[lut_1043_select];
    
    generate
    if ( USE_REG ) begin : ff_1043
        reg   lut_1043_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1043_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1043_ff <= lut_1043_out;
            end
        end
        
        assign out_data[1043] = lut_1043_ff;
    end
    else begin : no_ff_1043
        assign out_data[1043] = lut_1043_out;
    end
    endgenerate
    
    
    
    // LUT : 1044
    wire [63:0] lut_1044_table = 64'b0000111100001100111111111100111000001111000011110000111100001111;
    wire [5:0] lut_1044_select = {
                             in_data[487],
                             in_data[388],
                             in_data[770],
                             in_data[434],
                             in_data[640],
                             in_data[31]};
    
    wire lut_1044_out = lut_1044_table[lut_1044_select];
    
    generate
    if ( USE_REG ) begin : ff_1044
        reg   lut_1044_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1044_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1044_ff <= lut_1044_out;
            end
        end
        
        assign out_data[1044] = lut_1044_ff;
    end
    else begin : no_ff_1044
        assign out_data[1044] = lut_1044_out;
    end
    endgenerate
    
    
    
    // LUT : 1045
    wire [63:0] lut_1045_table = 64'b0000000011111111001000001111111100000000011101110000000011111111;
    wire [5:0] lut_1045_select = {
                             in_data[751],
                             in_data[114],
                             in_data[458],
                             in_data[16],
                             in_data[752],
                             in_data[60]};
    
    wire lut_1045_out = lut_1045_table[lut_1045_select];
    
    generate
    if ( USE_REG ) begin : ff_1045
        reg   lut_1045_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1045_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1045_ff <= lut_1045_out;
            end
        end
        
        assign out_data[1045] = lut_1045_ff;
    end
    else begin : no_ff_1045
        assign out_data[1045] = lut_1045_out;
    end
    endgenerate
    
    
    
    // LUT : 1046
    wire [63:0] lut_1046_table = 64'b0000000000000000000000000000000000000000000000001111111110111111;
    wire [5:0] lut_1046_select = {
                             in_data[678],
                             in_data[621],
                             in_data[531],
                             in_data[167],
                             in_data[233],
                             in_data[11]};
    
    wire lut_1046_out = lut_1046_table[lut_1046_select];
    
    generate
    if ( USE_REG ) begin : ff_1046
        reg   lut_1046_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1046_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1046_ff <= lut_1046_out;
            end
        end
        
        assign out_data[1046] = lut_1046_ff;
    end
    else begin : no_ff_1046
        assign out_data[1046] = lut_1046_out;
    end
    endgenerate
    
    
    
    // LUT : 1047
    wire [63:0] lut_1047_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1047_select = {
                             in_data[164],
                             in_data[206],
                             in_data[33],
                             in_data[310],
                             in_data[427],
                             in_data[36]};
    
    wire lut_1047_out = lut_1047_table[lut_1047_select];
    
    generate
    if ( USE_REG ) begin : ff_1047
        reg   lut_1047_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1047_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1047_ff <= lut_1047_out;
            end
        end
        
        assign out_data[1047] = lut_1047_ff;
    end
    else begin : no_ff_1047
        assign out_data[1047] = lut_1047_out;
    end
    endgenerate
    
    
    
    // LUT : 1048
    wire [63:0] lut_1048_table = 64'b0000111100001111000000000000111100001111000011110000000000001111;
    wire [5:0] lut_1048_select = {
                             in_data[9],
                             in_data[293],
                             in_data[556],
                             in_data[459],
                             in_data[725],
                             in_data[753]};
    
    wire lut_1048_out = lut_1048_table[lut_1048_select];
    
    generate
    if ( USE_REG ) begin : ff_1048
        reg   lut_1048_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1048_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1048_ff <= lut_1048_out;
            end
        end
        
        assign out_data[1048] = lut_1048_ff;
    end
    else begin : no_ff_1048
        assign out_data[1048] = lut_1048_out;
    end
    endgenerate
    
    
    
    // LUT : 1049
    wire [63:0] lut_1049_table = 64'b0011001100000000001100110000100000110011000000000011001110001000;
    wire [5:0] lut_1049_select = {
                             in_data[109],
                             in_data[693],
                             in_data[515],
                             in_data[35],
                             in_data[325],
                             in_data[598]};
    
    wire lut_1049_out = lut_1049_table[lut_1049_select];
    
    generate
    if ( USE_REG ) begin : ff_1049
        reg   lut_1049_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1049_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1049_ff <= lut_1049_out;
            end
        end
        
        assign out_data[1049] = lut_1049_ff;
    end
    else begin : no_ff_1049
        assign out_data[1049] = lut_1049_out;
    end
    endgenerate
    
    
    
    // LUT : 1050
    wire [63:0] lut_1050_table = 64'b1111111111001100111111111100110011101111110011001111110111001100;
    wire [5:0] lut_1050_select = {
                             in_data[334],
                             in_data[26],
                             in_data[157],
                             in_data[762],
                             in_data[629],
                             in_data[757]};
    
    wire lut_1050_out = lut_1050_table[lut_1050_select];
    
    generate
    if ( USE_REG ) begin : ff_1050
        reg   lut_1050_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1050_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1050_ff <= lut_1050_out;
            end
        end
        
        assign out_data[1050] = lut_1050_ff;
    end
    else begin : no_ff_1050
        assign out_data[1050] = lut_1050_out;
    end
    endgenerate
    
    
    
    // LUT : 1051
    wire [63:0] lut_1051_table = 64'b1111101111111011111110111111101111111011111110101111101011111010;
    wire [5:0] lut_1051_select = {
                             in_data[728],
                             in_data[727],
                             in_data[84],
                             in_data[744],
                             in_data[135],
                             in_data[592]};
    
    wire lut_1051_out = lut_1051_table[lut_1051_select];
    
    generate
    if ( USE_REG ) begin : ff_1051
        reg   lut_1051_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1051_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1051_ff <= lut_1051_out;
            end
        end
        
        assign out_data[1051] = lut_1051_ff;
    end
    else begin : no_ff_1051
        assign out_data[1051] = lut_1051_out;
    end
    endgenerate
    
    
    
    // LUT : 1052
    wire [63:0] lut_1052_table = 64'b1010101010101010111011101010111010101010101010101010111010101110;
    wire [5:0] lut_1052_select = {
                             in_data[738],
                             in_data[358],
                             in_data[572],
                             in_data[285],
                             in_data[511],
                             in_data[322]};
    
    wire lut_1052_out = lut_1052_table[lut_1052_select];
    
    generate
    if ( USE_REG ) begin : ff_1052
        reg   lut_1052_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1052_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1052_ff <= lut_1052_out;
            end
        end
        
        assign out_data[1052] = lut_1052_ff;
    end
    else begin : no_ff_1052
        assign out_data[1052] = lut_1052_out;
    end
    endgenerate
    
    
    
    // LUT : 1053
    wire [63:0] lut_1053_table = 64'b1111111111111111111111011101110111111111111111110101010101010100;
    wire [5:0] lut_1053_select = {
                             in_data[349],
                             in_data[158],
                             in_data[100],
                             in_data[473],
                             in_data[123],
                             in_data[658]};
    
    wire lut_1053_out = lut_1053_table[lut_1053_select];
    
    generate
    if ( USE_REG ) begin : ff_1053
        reg   lut_1053_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1053_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1053_ff <= lut_1053_out;
            end
        end
        
        assign out_data[1053] = lut_1053_ff;
    end
    else begin : no_ff_1053
        assign out_data[1053] = lut_1053_out;
    end
    endgenerate
    
    
    
    // LUT : 1054
    wire [63:0] lut_1054_table = 64'b1100111111001111111111111111111100001111000011110000011100000011;
    wire [5:0] lut_1054_select = {
                             in_data[568],
                             in_data[626],
                             in_data[674],
                             in_data[378],
                             in_data[635],
                             in_data[37]};
    
    wire lut_1054_out = lut_1054_table[lut_1054_select];
    
    generate
    if ( USE_REG ) begin : ff_1054
        reg   lut_1054_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1054_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1054_ff <= lut_1054_out;
            end
        end
        
        assign out_data[1054] = lut_1054_ff;
    end
    else begin : no_ff_1054
        assign out_data[1054] = lut_1054_out;
    end
    endgenerate
    
    
    
    // LUT : 1055
    wire [63:0] lut_1055_table = 64'b0011001100110000001100110011000000001111001111110000111100111111;
    wire [5:0] lut_1055_select = {
                             in_data[545],
                             in_data[182],
                             in_data[659],
                             in_data[576],
                             in_data[177],
                             in_data[774]};
    
    wire lut_1055_out = lut_1055_table[lut_1055_select];
    
    generate
    if ( USE_REG ) begin : ff_1055
        reg   lut_1055_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1055_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1055_ff <= lut_1055_out;
            end
        end
        
        assign out_data[1055] = lut_1055_ff;
    end
    else begin : no_ff_1055
        assign out_data[1055] = lut_1055_out;
    end
    endgenerate
    
    
    
    // LUT : 1056
    wire [63:0] lut_1056_table = 64'b0101010111010101010101001101110001010101111111010101010011011100;
    wire [5:0] lut_1056_select = {
                             in_data[506],
                             in_data[263],
                             in_data[105],
                             in_data[741],
                             in_data[318],
                             in_data[521]};
    
    wire lut_1056_out = lut_1056_table[lut_1056_select];
    
    generate
    if ( USE_REG ) begin : ff_1056
        reg   lut_1056_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1056_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1056_ff <= lut_1056_out;
            end
        end
        
        assign out_data[1056] = lut_1056_ff;
    end
    else begin : no_ff_1056
        assign out_data[1056] = lut_1056_out;
    end
    endgenerate
    
    
    
    // LUT : 1057
    wire [63:0] lut_1057_table = 64'b1111111111111111010100000101000011111111111111110101000001010000;
    wire [5:0] lut_1057_select = {
                             in_data[50],
                             in_data[552],
                             in_data[479],
                             in_data[429],
                             in_data[559],
                             in_data[265]};
    
    wire lut_1057_out = lut_1057_table[lut_1057_select];
    
    generate
    if ( USE_REG ) begin : ff_1057
        reg   lut_1057_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1057_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1057_ff <= lut_1057_out;
            end
        end
        
        assign out_data[1057] = lut_1057_ff;
    end
    else begin : no_ff_1057
        assign out_data[1057] = lut_1057_out;
    end
    endgenerate
    
    
    
    // LUT : 1058
    wire [63:0] lut_1058_table = 64'b1011111111111111101111111011111100111011101111110010001100100011;
    wire [5:0] lut_1058_select = {
                             in_data[636],
                             in_data[298],
                             in_data[430],
                             in_data[343],
                             in_data[401],
                             in_data[648]};
    
    wire lut_1058_out = lut_1058_table[lut_1058_select];
    
    generate
    if ( USE_REG ) begin : ff_1058
        reg   lut_1058_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1058_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1058_ff <= lut_1058_out;
            end
        end
        
        assign out_data[1058] = lut_1058_ff;
    end
    else begin : no_ff_1058
        assign out_data[1058] = lut_1058_out;
    end
    endgenerate
    
    
    
    // LUT : 1059
    wire [63:0] lut_1059_table = 64'b1111111100000101000010100000000011111111111111111111111101011111;
    wire [5:0] lut_1059_select = {
                             in_data[426],
                             in_data[582],
                             in_data[126],
                             in_data[357],
                             in_data[361],
                             in_data[300]};
    
    wire lut_1059_out = lut_1059_table[lut_1059_select];
    
    generate
    if ( USE_REG ) begin : ff_1059
        reg   lut_1059_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1059_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1059_ff <= lut_1059_out;
            end
        end
        
        assign out_data[1059] = lut_1059_ff;
    end
    else begin : no_ff_1059
        assign out_data[1059] = lut_1059_out;
    end
    endgenerate
    
    
    
    // LUT : 1060
    wire [63:0] lut_1060_table = 64'b0000000010101010000000001110101000000000101110100000000011111010;
    wire [5:0] lut_1060_select = {
                             in_data[24],
                             in_data[644],
                             in_data[236],
                             in_data[188],
                             in_data[391],
                             in_data[323]};
    
    wire lut_1060_out = lut_1060_table[lut_1060_select];
    
    generate
    if ( USE_REG ) begin : ff_1060
        reg   lut_1060_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1060_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1060_ff <= lut_1060_out;
            end
        end
        
        assign out_data[1060] = lut_1060_ff;
    end
    else begin : no_ff_1060
        assign out_data[1060] = lut_1060_out;
    end
    endgenerate
    
    
    
    // LUT : 1061
    wire [63:0] lut_1061_table = 64'b0000000000000000000010100000101010101010101010101010101010101010;
    wire [5:0] lut_1061_select = {
                             in_data[212],
                             in_data[416],
                             in_data[394],
                             in_data[424],
                             in_data[138],
                             in_data[516]};
    
    wire lut_1061_out = lut_1061_table[lut_1061_select];
    
    generate
    if ( USE_REG ) begin : ff_1061
        reg   lut_1061_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1061_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1061_ff <= lut_1061_out;
            end
        end
        
        assign out_data[1061] = lut_1061_ff;
    end
    else begin : no_ff_1061
        assign out_data[1061] = lut_1061_out;
    end
    endgenerate
    
    
    
    // LUT : 1062
    wire [63:0] lut_1062_table = 64'b1100110011001111000000000000000010000000000011110000000000000011;
    wire [5:0] lut_1062_select = {
                             in_data[716],
                             in_data[232],
                             in_data[289],
                             in_data[315],
                             in_data[690],
                             in_data[393]};
    
    wire lut_1062_out = lut_1062_table[lut_1062_select];
    
    generate
    if ( USE_REG ) begin : ff_1062
        reg   lut_1062_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1062_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1062_ff <= lut_1062_out;
            end
        end
        
        assign out_data[1062] = lut_1062_ff;
    end
    else begin : no_ff_1062
        assign out_data[1062] = lut_1062_out;
    end
    endgenerate
    
    
    
    // LUT : 1063
    wire [63:0] lut_1063_table = 64'b0101010101010101011101110100010001110111010101010111010100000000;
    wire [5:0] lut_1063_select = {
                             in_data[599],
                             in_data[383],
                             in_data[594],
                             in_data[88],
                             in_data[202],
                             in_data[347]};
    
    wire lut_1063_out = lut_1063_table[lut_1063_select];
    
    generate
    if ( USE_REG ) begin : ff_1063
        reg   lut_1063_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1063_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1063_ff <= lut_1063_out;
            end
        end
        
        assign out_data[1063] = lut_1063_ff;
    end
    else begin : no_ff_1063
        assign out_data[1063] = lut_1063_out;
    end
    endgenerate
    
    
    
    // LUT : 1064
    wire [63:0] lut_1064_table = 64'b0000101110000011001010111011101100001011100100111011101110111011;
    wire [5:0] lut_1064_select = {
                             in_data[63],
                             in_data[775],
                             in_data[269],
                             in_data[297],
                             in_data[351],
                             in_data[715]};
    
    wire lut_1064_out = lut_1064_table[lut_1064_select];
    
    generate
    if ( USE_REG ) begin : ff_1064
        reg   lut_1064_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1064_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1064_ff <= lut_1064_out;
            end
        end
        
        assign out_data[1064] = lut_1064_ff;
    end
    else begin : no_ff_1064
        assign out_data[1064] = lut_1064_out;
    end
    endgenerate
    
    
    
    // LUT : 1065
    wire [63:0] lut_1065_table = 64'b0100010011010101110000001111010011001100110111011101010011110101;
    wire [5:0] lut_1065_select = {
                             in_data[367],
                             in_data[550],
                             in_data[375],
                             in_data[132],
                             in_data[121],
                             in_data[101]};
    
    wire lut_1065_out = lut_1065_table[lut_1065_select];
    
    generate
    if ( USE_REG ) begin : ff_1065
        reg   lut_1065_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1065_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1065_ff <= lut_1065_out;
            end
        end
        
        assign out_data[1065] = lut_1065_ff;
    end
    else begin : no_ff_1065
        assign out_data[1065] = lut_1065_out;
    end
    endgenerate
    
    
    
    // LUT : 1066
    wire [63:0] lut_1066_table = 64'b1111001011111000111100001111000011010000111110001101000011110000;
    wire [5:0] lut_1066_select = {
                             in_data[483],
                             in_data[591],
                             in_data[551],
                             in_data[410],
                             in_data[163],
                             in_data[523]};
    
    wire lut_1066_out = lut_1066_table[lut_1066_select];
    
    generate
    if ( USE_REG ) begin : ff_1066
        reg   lut_1066_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1066_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1066_ff <= lut_1066_out;
            end
        end
        
        assign out_data[1066] = lut_1066_ff;
    end
    else begin : no_ff_1066
        assign out_data[1066] = lut_1066_out;
    end
    endgenerate
    
    
    
    // LUT : 1067
    wire [63:0] lut_1067_table = 64'b1100110001001100110011001000110011111111000000001111111100000000;
    wire [5:0] lut_1067_select = {
                             in_data[436],
                             in_data[166],
                             in_data[352],
                             in_data[477],
                             in_data[524],
                             in_data[144]};
    
    wire lut_1067_out = lut_1067_table[lut_1067_select];
    
    generate
    if ( USE_REG ) begin : ff_1067
        reg   lut_1067_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1067_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1067_ff <= lut_1067_out;
            end
        end
        
        assign out_data[1067] = lut_1067_ff;
    end
    else begin : no_ff_1067
        assign out_data[1067] = lut_1067_out;
    end
    endgenerate
    
    
    
    // LUT : 1068
    wire [63:0] lut_1068_table = 64'b0011001100000011001100110000001100110011000000110011001100000011;
    wire [5:0] lut_1068_select = {
                             in_data[15],
                             in_data[22],
                             in_data[340],
                             in_data[65],
                             in_data[497],
                             in_data[57]};
    
    wire lut_1068_out = lut_1068_table[lut_1068_select];
    
    generate
    if ( USE_REG ) begin : ff_1068
        reg   lut_1068_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1068_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1068_ff <= lut_1068_out;
            end
        end
        
        assign out_data[1068] = lut_1068_ff;
    end
    else begin : no_ff_1068
        assign out_data[1068] = lut_1068_out;
    end
    endgenerate
    
    
    
    // LUT : 1069
    wire [63:0] lut_1069_table = 64'b1111111111111111111111110000000011111111111111111111111110001000;
    wire [5:0] lut_1069_select = {
                             in_data[480],
                             in_data[597],
                             in_data[529],
                             in_data[45],
                             in_data[633],
                             in_data[279]};
    
    wire lut_1069_out = lut_1069_table[lut_1069_select];
    
    generate
    if ( USE_REG ) begin : ff_1069
        reg   lut_1069_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1069_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1069_ff <= lut_1069_out;
            end
        end
        
        assign out_data[1069] = lut_1069_ff;
    end
    else begin : no_ff_1069
        assign out_data[1069] = lut_1069_out;
    end
    endgenerate
    
    
    
    // LUT : 1070
    wire [63:0] lut_1070_table = 64'b1111101010111010111111111111111111111010101110101111111111111110;
    wire [5:0] lut_1070_select = {
                             in_data[764],
                             in_data[152],
                             in_data[714],
                             in_data[739],
                             in_data[631],
                             in_data[217]};
    
    wire lut_1070_out = lut_1070_table[lut_1070_select];
    
    generate
    if ( USE_REG ) begin : ff_1070
        reg   lut_1070_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1070_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1070_ff <= lut_1070_out;
            end
        end
        
        assign out_data[1070] = lut_1070_ff;
    end
    else begin : no_ff_1070
        assign out_data[1070] = lut_1070_out;
    end
    endgenerate
    
    
    
    // LUT : 1071
    wire [63:0] lut_1071_table = 64'b0011111110111111001100110011001100110011001100110000000000000000;
    wire [5:0] lut_1071_select = {
                             in_data[535],
                             in_data[291],
                             in_data[478],
                             in_data[585],
                             in_data[266],
                             in_data[362]};
    
    wire lut_1071_out = lut_1071_table[lut_1071_select];
    
    generate
    if ( USE_REG ) begin : ff_1071
        reg   lut_1071_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1071_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1071_ff <= lut_1071_out;
            end
        end
        
        assign out_data[1071] = lut_1071_ff;
    end
    else begin : no_ff_1071
        assign out_data[1071] = lut_1071_out;
    end
    endgenerate
    
    
    
    // LUT : 1072
    wire [63:0] lut_1072_table = 64'b0000000000000000111111111111111100000000000000001111010011110101;
    wire [5:0] lut_1072_select = {
                             in_data[264],
                             in_data[160],
                             in_data[505],
                             in_data[717],
                             in_data[729],
                             in_data[321]};
    
    wire lut_1072_out = lut_1072_table[lut_1072_select];
    
    generate
    if ( USE_REG ) begin : ff_1072
        reg   lut_1072_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1072_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1072_ff <= lut_1072_out;
            end
        end
        
        assign out_data[1072] = lut_1072_ff;
    end
    else begin : no_ff_1072
        assign out_data[1072] = lut_1072_out;
    end
    endgenerate
    
    
    
    // LUT : 1073
    wire [63:0] lut_1073_table = 64'b0000000000000000000000000000000000000000101111110000000011111111;
    wire [5:0] lut_1073_select = {
                             in_data[417],
                             in_data[779],
                             in_data[204],
                             in_data[694],
                             in_data[773],
                             in_data[197]};
    
    wire lut_1073_out = lut_1073_table[lut_1073_select];
    
    generate
    if ( USE_REG ) begin : ff_1073
        reg   lut_1073_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1073_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1073_ff <= lut_1073_out;
            end
        end
        
        assign out_data[1073] = lut_1073_ff;
    end
    else begin : no_ff_1073
        assign out_data[1073] = lut_1073_out;
    end
    endgenerate
    
    
    
    // LUT : 1074
    wire [63:0] lut_1074_table = 64'b0000100000000000000000001000100011101110111011101110111011101110;
    wire [5:0] lut_1074_select = {
                             in_data[294],
                             in_data[85],
                             in_data[143],
                             in_data[395],
                             in_data[745],
                             in_data[382]};
    
    wire lut_1074_out = lut_1074_table[lut_1074_select];
    
    generate
    if ( USE_REG ) begin : ff_1074
        reg   lut_1074_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1074_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1074_ff <= lut_1074_out;
            end
        end
        
        assign out_data[1074] = lut_1074_ff;
    end
    else begin : no_ff_1074
        assign out_data[1074] = lut_1074_out;
    end
    endgenerate
    
    
    
    // LUT : 1075
    wire [63:0] lut_1075_table = 64'b0000000000000000111111111111000011000000000000001111111111110000;
    wire [5:0] lut_1075_select = {
                             in_data[32],
                             in_data[368],
                             in_data[610],
                             in_data[208],
                             in_data[514],
                             in_data[783]};
    
    wire lut_1075_out = lut_1075_table[lut_1075_select];
    
    generate
    if ( USE_REG ) begin : ff_1075
        reg   lut_1075_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1075_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1075_ff <= lut_1075_out;
            end
        end
        
        assign out_data[1075] = lut_1075_ff;
    end
    else begin : no_ff_1075
        assign out_data[1075] = lut_1075_out;
    end
    endgenerate
    
    
    
    // LUT : 1076
    wire [63:0] lut_1076_table = 64'b1100000011001100110011001100110000000000000000001111111111001100;
    wire [5:0] lut_1076_select = {
                             in_data[178],
                             in_data[580],
                             in_data[324],
                             in_data[92],
                             in_data[379],
                             in_data[227]};
    
    wire lut_1076_out = lut_1076_table[lut_1076_select];
    
    generate
    if ( USE_REG ) begin : ff_1076
        reg   lut_1076_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1076_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1076_ff <= lut_1076_out;
            end
        end
        
        assign out_data[1076] = lut_1076_ff;
    end
    else begin : no_ff_1076
        assign out_data[1076] = lut_1076_out;
    end
    endgenerate
    
    
    
    // LUT : 1077
    wire [63:0] lut_1077_table = 64'b1111111111001100111111111100110011001100110011001100110011001100;
    wire [5:0] lut_1077_select = {
                             in_data[467],
                             in_data[19],
                             in_data[237],
                             in_data[339],
                             in_data[565],
                             in_data[113]};
    
    wire lut_1077_out = lut_1077_table[lut_1077_select];
    
    generate
    if ( USE_REG ) begin : ff_1077
        reg   lut_1077_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1077_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1077_ff <= lut_1077_out;
            end
        end
        
        assign out_data[1077] = lut_1077_ff;
    end
    else begin : no_ff_1077
        assign out_data[1077] = lut_1077_out;
    end
    endgenerate
    
    
    
    // LUT : 1078
    wire [63:0] lut_1078_table = 64'b0000110100001101000011010000110100001100000011010000110100001101;
    wire [5:0] lut_1078_select = {
                             in_data[127],
                             in_data[116],
                             in_data[137],
                             in_data[488],
                             in_data[181],
                             in_data[498]};
    
    wire lut_1078_out = lut_1078_table[lut_1078_select];
    
    generate
    if ( USE_REG ) begin : ff_1078
        reg   lut_1078_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1078_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1078_ff <= lut_1078_out;
            end
        end
        
        assign out_data[1078] = lut_1078_ff;
    end
    else begin : no_ff_1078
        assign out_data[1078] = lut_1078_out;
    end
    endgenerate
    
    
    
    // LUT : 1079
    wire [63:0] lut_1079_table = 64'b1010101011111111111111111111111100000000101011100000000010101010;
    wire [5:0] lut_1079_select = {
                             in_data[218],
                             in_data[268],
                             in_data[247],
                             in_data[670],
                             in_data[418],
                             in_data[244]};
    
    wire lut_1079_out = lut_1079_table[lut_1079_select];
    
    generate
    if ( USE_REG ) begin : ff_1079
        reg   lut_1079_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1079_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1079_ff <= lut_1079_out;
            end
        end
        
        assign out_data[1079] = lut_1079_ff;
    end
    else begin : no_ff_1079
        assign out_data[1079] = lut_1079_out;
    end
    endgenerate
    
    
    
    // LUT : 1080
    wire [63:0] lut_1080_table = 64'b0000111111111111101011111111111110101111101011111010101010101010;
    wire [5:0] lut_1080_select = {
                             in_data[441],
                             in_data[494],
                             in_data[187],
                             in_data[464],
                             in_data[43],
                             in_data[712]};
    
    wire lut_1080_out = lut_1080_table[lut_1080_select];
    
    generate
    if ( USE_REG ) begin : ff_1080
        reg   lut_1080_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1080_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1080_ff <= lut_1080_out;
            end
        end
        
        assign out_data[1080] = lut_1080_ff;
    end
    else begin : no_ff_1080
        assign out_data[1080] = lut_1080_out;
    end
    endgenerate
    
    
    
    // LUT : 1081
    wire [63:0] lut_1081_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_1081_select = {
                             in_data[442],
                             in_data[222],
                             in_data[21],
                             in_data[642],
                             in_data[12],
                             in_data[34]};
    
    wire lut_1081_out = lut_1081_table[lut_1081_select];
    
    generate
    if ( USE_REG ) begin : ff_1081
        reg   lut_1081_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1081_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1081_ff <= lut_1081_out;
            end
        end
        
        assign out_data[1081] = lut_1081_ff;
    end
    else begin : no_ff_1081
        assign out_data[1081] = lut_1081_out;
    end
    endgenerate
    
    
    
    // LUT : 1082
    wire [63:0] lut_1082_table = 64'b1111110011111111111111111111111111110000111100001111000011110000;
    wire [5:0] lut_1082_select = {
                             in_data[713],
                             in_data[680],
                             in_data[40],
                             in_data[398],
                             in_data[443],
                             in_data[223]};
    
    wire lut_1082_out = lut_1082_table[lut_1082_select];
    
    generate
    if ( USE_REG ) begin : ff_1082
        reg   lut_1082_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1082_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1082_ff <= lut_1082_out;
            end
        end
        
        assign out_data[1082] = lut_1082_ff;
    end
    else begin : no_ff_1082
        assign out_data[1082] = lut_1082_out;
    end
    endgenerate
    
    
    
    // LUT : 1083
    wire [63:0] lut_1083_table = 64'b0000000000000000000100110001001100000100000001000001011100010111;
    wire [5:0] lut_1083_select = {
                             in_data[161],
                             in_data[484],
                             in_data[449],
                             in_data[74],
                             in_data[453],
                             in_data[387]};
    
    wire lut_1083_out = lut_1083_table[lut_1083_select];
    
    generate
    if ( USE_REG ) begin : ff_1083
        reg   lut_1083_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1083_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1083_ff <= lut_1083_out;
            end
        end
        
        assign out_data[1083] = lut_1083_ff;
    end
    else begin : no_ff_1083
        assign out_data[1083] = lut_1083_out;
    end
    endgenerate
    
    
    
    // LUT : 1084
    wire [63:0] lut_1084_table = 64'b0000010111111111000111111111111100000000011100000000000011110000;
    wire [5:0] lut_1084_select = {
                             in_data[639],
                             in_data[304],
                             in_data[596],
                             in_data[373],
                             in_data[765],
                             in_data[201]};
    
    wire lut_1084_out = lut_1084_table[lut_1084_select];
    
    generate
    if ( USE_REG ) begin : ff_1084
        reg   lut_1084_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1084_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1084_ff <= lut_1084_out;
            end
        end
        
        assign out_data[1084] = lut_1084_ff;
    end
    else begin : no_ff_1084
        assign out_data[1084] = lut_1084_out;
    end
    endgenerate
    
    
    
    // LUT : 1085
    wire [63:0] lut_1085_table = 64'b0010111110101111101011111010111110101111101011111010111110101111;
    wire [5:0] lut_1085_select = {
                             in_data[731],
                             in_data[111],
                             in_data[59],
                             in_data[435],
                             in_data[557],
                             in_data[246]};
    
    wire lut_1085_out = lut_1085_table[lut_1085_select];
    
    generate
    if ( USE_REG ) begin : ff_1085
        reg   lut_1085_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1085_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1085_ff <= lut_1085_out;
            end
        end
        
        assign out_data[1085] = lut_1085_ff;
    end
    else begin : no_ff_1085
        assign out_data[1085] = lut_1085_out;
    end
    endgenerate
    
    
    
    // LUT : 1086
    wire [63:0] lut_1086_table = 64'b1111111111111111000000001111111111111111111111110010101010101010;
    wire [5:0] lut_1086_select = {
                             in_data[369],
                             in_data[150],
                             in_data[260],
                             in_data[30],
                             in_data[140],
                             in_data[415]};
    
    wire lut_1086_out = lut_1086_table[lut_1086_select];
    
    generate
    if ( USE_REG ) begin : ff_1086
        reg   lut_1086_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1086_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1086_ff <= lut_1086_out;
            end
        end
        
        assign out_data[1086] = lut_1086_ff;
    end
    else begin : no_ff_1086
        assign out_data[1086] = lut_1086_out;
    end
    endgenerate
    
    
    
    // LUT : 1087
    wire [63:0] lut_1087_table = 64'b0111011101100110111111110110011001000100000000000101010101010101;
    wire [5:0] lut_1087_select = {
                             in_data[625],
                             in_data[312],
                             in_data[660],
                             in_data[56],
                             in_data[372],
                             in_data[437]};
    
    wire lut_1087_out = lut_1087_table[lut_1087_select];
    
    generate
    if ( USE_REG ) begin : ff_1087
        reg   lut_1087_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1087_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1087_ff <= lut_1087_out;
            end
        end
        
        assign out_data[1087] = lut_1087_ff;
    end
    else begin : no_ff_1087
        assign out_data[1087] = lut_1087_out;
    end
    endgenerate
    
    
    
    // LUT : 1088
    wire [63:0] lut_1088_table = 64'b0000000000000000000000100000101000000000000000000000001000001010;
    wire [5:0] lut_1088_select = {
                             in_data[78],
                             in_data[653],
                             in_data[170],
                             in_data[189],
                             in_data[507],
                             in_data[457]};
    
    wire lut_1088_out = lut_1088_table[lut_1088_select];
    
    generate
    if ( USE_REG ) begin : ff_1088
        reg   lut_1088_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1088_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1088_ff <= lut_1088_out;
            end
        end
        
        assign out_data[1088] = lut_1088_ff;
    end
    else begin : no_ff_1088
        assign out_data[1088] = lut_1088_out;
    end
    endgenerate
    
    
    
    // LUT : 1089
    wire [63:0] lut_1089_table = 64'b1111111111111111111111111100110011111111111111111111111111001110;
    wire [5:0] lut_1089_select = {
                             in_data[280],
                             in_data[452],
                             in_data[685],
                             in_data[41],
                             in_data[250],
                             in_data[419]};
    
    wire lut_1089_out = lut_1089_table[lut_1089_select];
    
    generate
    if ( USE_REG ) begin : ff_1089
        reg   lut_1089_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1089_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1089_ff <= lut_1089_out;
            end
        end
        
        assign out_data[1089] = lut_1089_ff;
    end
    else begin : no_ff_1089
        assign out_data[1089] = lut_1089_out;
    end
    endgenerate
    
    
    
    // LUT : 1090
    wire [63:0] lut_1090_table = 64'b1111111111111111101000001111101111111111111111111010000011111111;
    wire [5:0] lut_1090_select = {
                             in_data[760],
                             in_data[190],
                             in_data[210],
                             in_data[593],
                             in_data[673],
                             in_data[405]};
    
    wire lut_1090_out = lut_1090_table[lut_1090_select];
    
    generate
    if ( USE_REG ) begin : ff_1090
        reg   lut_1090_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1090_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1090_ff <= lut_1090_out;
            end
        end
        
        assign out_data[1090] = lut_1090_ff;
    end
    else begin : no_ff_1090
        assign out_data[1090] = lut_1090_out;
    end
    endgenerate
    
    
    
    // LUT : 1091
    wire [63:0] lut_1091_table = 64'b0011001100110000001100110011000000110011111100001111001111110011;
    wire [5:0] lut_1091_select = {
                             in_data[574],
                             in_data[68],
                             in_data[519],
                             in_data[691],
                             in_data[99],
                             in_data[561]};
    
    wire lut_1091_out = lut_1091_table[lut_1091_select];
    
    generate
    if ( USE_REG ) begin : ff_1091
        reg   lut_1091_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1091_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1091_ff <= lut_1091_out;
            end
        end
        
        assign out_data[1091] = lut_1091_ff;
    end
    else begin : no_ff_1091
        assign out_data[1091] = lut_1091_out;
    end
    endgenerate
    
    
    
    // LUT : 1092
    wire [63:0] lut_1092_table = 64'b0111011101010101010101010000000011110111010101010101010100000000;
    wire [5:0] lut_1092_select = {
                             in_data[38],
                             in_data[581],
                             in_data[721],
                             in_data[364],
                             in_data[749],
                             in_data[681]};
    
    wire lut_1092_out = lut_1092_table[lut_1092_select];
    
    generate
    if ( USE_REG ) begin : ff_1092
        reg   lut_1092_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1092_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1092_ff <= lut_1092_out;
            end
        end
        
        assign out_data[1092] = lut_1092_ff;
    end
    else begin : no_ff_1092
        assign out_data[1092] = lut_1092_out;
    end
    endgenerate
    
    
    
    // LUT : 1093
    wire [63:0] lut_1093_table = 64'b0100010011111111010001001101110101000100111111110000000011011101;
    wire [5:0] lut_1093_select = {
                             in_data[615],
                             in_data[696],
                             in_data[440],
                             in_data[474],
                             in_data[97],
                             in_data[722]};
    
    wire lut_1093_out = lut_1093_table[lut_1093_select];
    
    generate
    if ( USE_REG ) begin : ff_1093
        reg   lut_1093_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1093_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1093_ff <= lut_1093_out;
            end
        end
        
        assign out_data[1093] = lut_1093_ff;
    end
    else begin : no_ff_1093
        assign out_data[1093] = lut_1093_out;
    end
    endgenerate
    
    
    
    // LUT : 1094
    wire [63:0] lut_1094_table = 64'b0000000000010000000100010001000100000000000000000001000100010001;
    wire [5:0] lut_1094_select = {
                             in_data[643],
                             in_data[207],
                             in_data[62],
                             in_data[723],
                             in_data[611],
                             in_data[70]};
    
    wire lut_1094_out = lut_1094_table[lut_1094_select];
    
    generate
    if ( USE_REG ) begin : ff_1094
        reg   lut_1094_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1094_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1094_ff <= lut_1094_out;
            end
        end
        
        assign out_data[1094] = lut_1094_ff;
    end
    else begin : no_ff_1094
        assign out_data[1094] = lut_1094_out;
    end
    endgenerate
    
    
    
    // LUT : 1095
    wire [63:0] lut_1095_table = 64'b1111111110101111111011111010101111111111101011111110111110101011;
    wire [5:0] lut_1095_select = {
                             in_data[6],
                             in_data[679],
                             in_data[286],
                             in_data[214],
                             in_data[495],
                             in_data[595]};
    
    wire lut_1095_out = lut_1095_table[lut_1095_select];
    
    generate
    if ( USE_REG ) begin : ff_1095
        reg   lut_1095_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1095_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1095_ff <= lut_1095_out;
            end
        end
        
        assign out_data[1095] = lut_1095_ff;
    end
    else begin : no_ff_1095
        assign out_data[1095] = lut_1095_out;
    end
    endgenerate
    
    
    
    // LUT : 1096
    wire [63:0] lut_1096_table = 64'b0000000000000000101011101010101000001100000001001111111111111111;
    wire [5:0] lut_1096_select = {
                             in_data[159],
                             in_data[413],
                             in_data[502],
                             in_data[632],
                             in_data[200],
                             in_data[354]};
    
    wire lut_1096_out = lut_1096_table[lut_1096_select];
    
    generate
    if ( USE_REG ) begin : ff_1096
        reg   lut_1096_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1096_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1096_ff <= lut_1096_out;
            end
        end
        
        assign out_data[1096] = lut_1096_ff;
    end
    else begin : no_ff_1096
        assign out_data[1096] = lut_1096_out;
    end
    endgenerate
    
    
    
    // LUT : 1097
    wire [63:0] lut_1097_table = 64'b1010111011101111101011111110111100001000100010100000100010001110;
    wire [5:0] lut_1097_select = {
                             in_data[290],
                             in_data[284],
                             in_data[95],
                             in_data[91],
                             in_data[245],
                             in_data[329]};
    
    wire lut_1097_out = lut_1097_table[lut_1097_select];
    
    generate
    if ( USE_REG ) begin : ff_1097
        reg   lut_1097_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1097_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1097_ff <= lut_1097_out;
            end
        end
        
        assign out_data[1097] = lut_1097_ff;
    end
    else begin : no_ff_1097
        assign out_data[1097] = lut_1097_out;
    end
    endgenerate
    
    
    
    // LUT : 1098
    wire [63:0] lut_1098_table = 64'b0000111100001100000011100000110011001111111111110100111111111111;
    wire [5:0] lut_1098_select = {
                             in_data[411],
                             in_data[776],
                             in_data[664],
                             in_data[605],
                             in_data[708],
                             in_data[184]};
    
    wire lut_1098_out = lut_1098_table[lut_1098_select];
    
    generate
    if ( USE_REG ) begin : ff_1098
        reg   lut_1098_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1098_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1098_ff <= lut_1098_out;
            end
        end
        
        assign out_data[1098] = lut_1098_ff;
    end
    else begin : no_ff_1098
        assign out_data[1098] = lut_1098_out;
    end
    endgenerate
    
    
    
    // LUT : 1099
    wire [63:0] lut_1099_table = 64'b1100111011001111110010001100110011001111110011111100010011001100;
    wire [5:0] lut_1099_select = {
                             in_data[684],
                             in_data[692],
                             in_data[433],
                             in_data[439],
                             in_data[183],
                             in_data[601]};
    
    wire lut_1099_out = lut_1099_table[lut_1099_select];
    
    generate
    if ( USE_REG ) begin : ff_1099
        reg   lut_1099_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1099_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1099_ff <= lut_1099_out;
            end
        end
        
        assign out_data[1099] = lut_1099_ff;
    end
    else begin : no_ff_1099
        assign out_data[1099] = lut_1099_out;
    end
    endgenerate
    
    
    
    // LUT : 1100
    wire [63:0] lut_1100_table = 64'b0000000000000000000000000000000011001100110011001100110011001100;
    wire [5:0] lut_1100_select = {
                             in_data[331],
                             in_data[44],
                             in_data[48],
                             in_data[650],
                             in_data[482],
                             in_data[700]};
    
    wire lut_1100_out = lut_1100_table[lut_1100_select];
    
    generate
    if ( USE_REG ) begin : ff_1100
        reg   lut_1100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1100_ff <= lut_1100_out;
            end
        end
        
        assign out_data[1100] = lut_1100_ff;
    end
    else begin : no_ff_1100
        assign out_data[1100] = lut_1100_out;
    end
    endgenerate
    
    
    
    // LUT : 1101
    wire [63:0] lut_1101_table = 64'b0011001100111011001100110011101100111011001110110011001100111011;
    wire [5:0] lut_1101_select = {
                             in_data[252],
                             in_data[709],
                             in_data[133],
                             in_data[462],
                             in_data[376],
                             in_data[128]};
    
    wire lut_1101_out = lut_1101_table[lut_1101_select];
    
    generate
    if ( USE_REG ) begin : ff_1101
        reg   lut_1101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1101_ff <= lut_1101_out;
            end
        end
        
        assign out_data[1101] = lut_1101_ff;
    end
    else begin : no_ff_1101
        assign out_data[1101] = lut_1101_out;
    end
    endgenerate
    
    
    
    // LUT : 1102
    wire [63:0] lut_1102_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_1102_select = {
                             in_data[371],
                             in_data[645],
                             in_data[274],
                             in_data[614],
                             in_data[667],
                             in_data[444]};
    
    wire lut_1102_out = lut_1102_table[lut_1102_select];
    
    generate
    if ( USE_REG ) begin : ff_1102
        reg   lut_1102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1102_ff <= lut_1102_out;
            end
        end
        
        assign out_data[1102] = lut_1102_ff;
    end
    else begin : no_ff_1102
        assign out_data[1102] = lut_1102_out;
    end
    endgenerate
    
    
    
    // LUT : 1103
    wire [63:0] lut_1103_table = 64'b0111111101111111000000000000100001111111011111110101100000011010;
    wire [5:0] lut_1103_select = {
                             in_data[10],
                             in_data[319],
                             in_data[569],
                             in_data[328],
                             in_data[104],
                             in_data[156]};
    
    wire lut_1103_out = lut_1103_table[lut_1103_select];
    
    generate
    if ( USE_REG ) begin : ff_1103
        reg   lut_1103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1103_ff <= lut_1103_out;
            end
        end
        
        assign out_data[1103] = lut_1103_ff;
    end
    else begin : no_ff_1103
        assign out_data[1103] = lut_1103_out;
    end
    endgenerate
    
    
    
    // LUT : 1104
    wire [63:0] lut_1104_table = 64'b1111111111111111101010111010101011111111111111110000000010000000;
    wire [5:0] lut_1104_select = {
                             in_data[93],
                             in_data[460],
                             in_data[534],
                             in_data[408],
                             in_data[558],
                             in_data[380]};
    
    wire lut_1104_out = lut_1104_table[lut_1104_select];
    
    generate
    if ( USE_REG ) begin : ff_1104
        reg   lut_1104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1104_ff <= lut_1104_out;
            end
        end
        
        assign out_data[1104] = lut_1104_ff;
    end
    else begin : no_ff_1104
        assign out_data[1104] = lut_1104_out;
    end
    endgenerate
    
    
    
    // LUT : 1105
    wire [63:0] lut_1105_table = 64'b0000111100001111111111111111111100001111000011111111111111111111;
    wire [5:0] lut_1105_select = {
                             in_data[771],
                             in_data[549],
                             in_data[384],
                             in_data[493],
                             in_data[49],
                             in_data[641]};
    
    wire lut_1105_out = lut_1105_table[lut_1105_select];
    
    generate
    if ( USE_REG ) begin : ff_1105
        reg   lut_1105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1105_ff <= lut_1105_out;
            end
        end
        
        assign out_data[1105] = lut_1105_ff;
    end
    else begin : no_ff_1105
        assign out_data[1105] = lut_1105_out;
    end
    endgenerate
    
    
    
    // LUT : 1106
    wire [63:0] lut_1106_table = 64'b0101111100001010010111110000101001011111000010100101111100001010;
    wire [5:0] lut_1106_select = {
                             in_data[25],
                             in_data[587],
                             in_data[657],
                             in_data[148],
                             in_data[29],
                             in_data[666]};
    
    wire lut_1106_out = lut_1106_table[lut_1106_select];
    
    generate
    if ( USE_REG ) begin : ff_1106
        reg   lut_1106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1106_ff <= lut_1106_out;
            end
        end
        
        assign out_data[1106] = lut_1106_ff;
    end
    else begin : no_ff_1106
        assign out_data[1106] = lut_1106_out;
    end
    endgenerate
    
    
    
    // LUT : 1107
    wire [63:0] lut_1107_table = 64'b0101110011011100110111001111111111011100110111001101110011111111;
    wire [5:0] lut_1107_select = {
                             in_data[47],
                             in_data[238],
                             in_data[768],
                             in_data[432],
                             in_data[663],
                             in_data[240]};
    
    wire lut_1107_out = lut_1107_table[lut_1107_select];
    
    generate
    if ( USE_REG ) begin : ff_1107
        reg   lut_1107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1107_ff <= lut_1107_out;
            end
        end
        
        assign out_data[1107] = lut_1107_ff;
    end
    else begin : no_ff_1107
        assign out_data[1107] = lut_1107_out;
    end
    endgenerate
    
    
    
    // LUT : 1108
    wire [63:0] lut_1108_table = 64'b0000000000000000000010110000101100000000000000000000111100001111;
    wire [5:0] lut_1108_select = {
                             in_data[704],
                             in_data[510],
                             in_data[589],
                             in_data[98],
                             in_data[147],
                             in_data[13]};
    
    wire lut_1108_out = lut_1108_table[lut_1108_select];
    
    generate
    if ( USE_REG ) begin : ff_1108
        reg   lut_1108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1108_ff <= lut_1108_out;
            end
        end
        
        assign out_data[1108] = lut_1108_ff;
    end
    else begin : no_ff_1108
        assign out_data[1108] = lut_1108_out;
    end
    endgenerate
    
    
    
    // LUT : 1109
    wire [63:0] lut_1109_table = 64'b1111111111111111001100110011001111111111111111110011001100110011;
    wire [5:0] lut_1109_select = {
                             in_data[763],
                             in_data[248],
                             in_data[527],
                             in_data[309],
                             in_data[512],
                             in_data[139]};
    
    wire lut_1109_out = lut_1109_table[lut_1109_select];
    
    generate
    if ( USE_REG ) begin : ff_1109
        reg   lut_1109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1109_ff <= lut_1109_out;
            end
        end
        
        assign out_data[1109] = lut_1109_ff;
    end
    else begin : no_ff_1109
        assign out_data[1109] = lut_1109_out;
    end
    endgenerate
    
    
    
    // LUT : 1110
    wire [63:0] lut_1110_table = 64'b1011101110111011001100110011001110110011101100110010001100110011;
    wire [5:0] lut_1110_select = {
                             in_data[651],
                             in_data[537],
                             in_data[754],
                             in_data[469],
                             in_data[153],
                             in_data[548]};
    
    wire lut_1110_out = lut_1110_table[lut_1110_select];
    
    generate
    if ( USE_REG ) begin : ff_1110
        reg   lut_1110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1110_ff <= lut_1110_out;
            end
        end
        
        assign out_data[1110] = lut_1110_ff;
    end
    else begin : no_ff_1110
        assign out_data[1110] = lut_1110_out;
    end
    endgenerate
    
    
    
    // LUT : 1111
    wire [63:0] lut_1111_table = 64'b1101110111011100010001000100010011011101110111010101010101010101;
    wire [5:0] lut_1111_select = {
                             in_data[149],
                             in_data[466],
                             in_data[737],
                             in_data[256],
                             in_data[314],
                             in_data[606]};
    
    wire lut_1111_out = lut_1111_table[lut_1111_select];
    
    generate
    if ( USE_REG ) begin : ff_1111
        reg   lut_1111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1111_ff <= lut_1111_out;
            end
        end
        
        assign out_data[1111] = lut_1111_ff;
    end
    else begin : no_ff_1111
        assign out_data[1111] = lut_1111_out;
    end
    endgenerate
    
    
    
    // LUT : 1112
    wire [63:0] lut_1112_table = 64'b1100111011101110000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1112_select = {
                             in_data[262],
                             in_data[131],
                             in_data[281],
                             in_data[778],
                             in_data[470],
                             in_data[54]};
    
    wire lut_1112_out = lut_1112_table[lut_1112_select];
    
    generate
    if ( USE_REG ) begin : ff_1112
        reg   lut_1112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1112_ff <= lut_1112_out;
            end
        end
        
        assign out_data[1112] = lut_1112_ff;
    end
    else begin : no_ff_1112
        assign out_data[1112] = lut_1112_out;
    end
    endgenerate
    
    
    
    // LUT : 1113
    wire [63:0] lut_1113_table = 64'b1111001100110011111100001111000011110011001100111110000011110101;
    wire [5:0] lut_1113_select = {
                             in_data[169],
                             in_data[216],
                             in_data[209],
                             in_data[688],
                             in_data[567],
                             in_data[81]};
    
    wire lut_1113_out = lut_1113_table[lut_1113_select];
    
    generate
    if ( USE_REG ) begin : ff_1113
        reg   lut_1113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1113_ff <= lut_1113_out;
            end
        end
        
        assign out_data[1113] = lut_1113_ff;
    end
    else begin : no_ff_1113
        assign out_data[1113] = lut_1113_out;
    end
    endgenerate
    
    
    
    // LUT : 1114
    wire [63:0] lut_1114_table = 64'b0101111100000101010111110000010001011111000001010101110100000000;
    wire [5:0] lut_1114_select = {
                             in_data[27],
                             in_data[0],
                             in_data[520],
                             in_data[303],
                             in_data[225],
                             in_data[235]};
    
    wire lut_1114_out = lut_1114_table[lut_1114_select];
    
    generate
    if ( USE_REG ) begin : ff_1114
        reg   lut_1114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1114_ff <= lut_1114_out;
            end
        end
        
        assign out_data[1114] = lut_1114_ff;
    end
    else begin : no_ff_1114
        assign out_data[1114] = lut_1114_out;
    end
    endgenerate
    
    
    
    // LUT : 1115
    wire [63:0] lut_1115_table = 64'b0000001100000111000000110001001100000011000001110000001100010011;
    wire [5:0] lut_1115_select = {
                             in_data[476],
                             in_data[547],
                             in_data[736],
                             in_data[627],
                             in_data[348],
                             in_data[277]};
    
    wire lut_1115_out = lut_1115_table[lut_1115_select];
    
    generate
    if ( USE_REG ) begin : ff_1115
        reg   lut_1115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1115_ff <= lut_1115_out;
            end
        end
        
        assign out_data[1115] = lut_1115_ff;
    end
    else begin : no_ff_1115
        assign out_data[1115] = lut_1115_out;
    end
    endgenerate
    
    
    
    // LUT : 1116
    wire [63:0] lut_1116_table = 64'b1111111101010101111111110101010101011111000000000101010101010000;
    wire [5:0] lut_1116_select = {
                             in_data[468],
                             in_data[518],
                             in_data[508],
                             in_data[342],
                             in_data[697],
                             in_data[463]};
    
    wire lut_1116_out = lut_1116_table[lut_1116_select];
    
    generate
    if ( USE_REG ) begin : ff_1116
        reg   lut_1116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1116_ff <= lut_1116_out;
            end
        end
        
        assign out_data[1116] = lut_1116_ff;
    end
    else begin : no_ff_1116
        assign out_data[1116] = lut_1116_out;
    end
    endgenerate
    
    
    
    // LUT : 1117
    wire [63:0] lut_1117_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_1117_select = {
                             in_data[226],
                             in_data[288],
                             in_data[399],
                             in_data[8],
                             in_data[726],
                             in_data[616]};
    
    wire lut_1117_out = lut_1117_table[lut_1117_select];
    
    generate
    if ( USE_REG ) begin : ff_1117
        reg   lut_1117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1117_ff <= lut_1117_out;
            end
        end
        
        assign out_data[1117] = lut_1117_ff;
    end
    else begin : no_ff_1117
        assign out_data[1117] = lut_1117_out;
    end
    endgenerate
    
    
    
    // LUT : 1118
    wire [63:0] lut_1118_table = 64'b1111111111111111111111111010000011111111111111111111111110100000;
    wire [5:0] lut_1118_select = {
                             in_data[392],
                             in_data[203],
                             in_data[179],
                             in_data[772],
                             in_data[513],
                             in_data[546]};
    
    wire lut_1118_out = lut_1118_table[lut_1118_select];
    
    generate
    if ( USE_REG ) begin : ff_1118
        reg   lut_1118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1118_ff <= lut_1118_out;
            end
        end
        
        assign out_data[1118] = lut_1118_ff;
    end
    else begin : no_ff_1118
        assign out_data[1118] = lut_1118_out;
    end
    endgenerate
    
    
    
    // LUT : 1119
    wire [63:0] lut_1119_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_1119_select = {
                             in_data[73],
                             in_data[486],
                             in_data[579],
                             in_data[702],
                             in_data[652],
                             in_data[261]};
    
    wire lut_1119_out = lut_1119_table[lut_1119_select];
    
    generate
    if ( USE_REG ) begin : ff_1119
        reg   lut_1119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1119_ff <= lut_1119_out;
            end
        end
        
        assign out_data[1119] = lut_1119_ff;
    end
    else begin : no_ff_1119
        assign out_data[1119] = lut_1119_out;
    end
    endgenerate
    
    
    
    // LUT : 1120
    wire [63:0] lut_1120_table = 64'b1111110111111111111111001111111111011100111111001100110011111100;
    wire [5:0] lut_1120_select = {
                             in_data[496],
                             in_data[82],
                             in_data[490],
                             in_data[528],
                             in_data[155],
                             in_data[112]};
    
    wire lut_1120_out = lut_1120_table[lut_1120_select];
    
    generate
    if ( USE_REG ) begin : ff_1120
        reg   lut_1120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1120_ff <= lut_1120_out;
            end
        end
        
        assign out_data[1120] = lut_1120_ff;
    end
    else begin : no_ff_1120
        assign out_data[1120] = lut_1120_out;
    end
    endgenerate
    
    
    
    // LUT : 1121
    wire [63:0] lut_1121_table = 64'b1111111111111111111111111111111100110011000000000011001000000000;
    wire [5:0] lut_1121_select = {
                             in_data[292],
                             in_data[46],
                             in_data[573],
                             in_data[390],
                             in_data[734],
                             in_data[421]};
    
    wire lut_1121_out = lut_1121_table[lut_1121_select];
    
    generate
    if ( USE_REG ) begin : ff_1121
        reg   lut_1121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1121_ff <= lut_1121_out;
            end
        end
        
        assign out_data[1121] = lut_1121_ff;
    end
    else begin : no_ff_1121
        assign out_data[1121] = lut_1121_out;
    end
    endgenerate
    
    
    
    // LUT : 1122
    wire [63:0] lut_1122_table = 64'b1111111111111111111111111111111111001100110011001111111111111111;
    wire [5:0] lut_1122_select = {
                             in_data[273],
                             in_data[239],
                             in_data[698],
                             in_data[646],
                             in_data[686],
                             in_data[316]};
    
    wire lut_1122_out = lut_1122_table[lut_1122_select];
    
    generate
    if ( USE_REG ) begin : ff_1122
        reg   lut_1122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1122_ff <= lut_1122_out;
            end
        end
        
        assign out_data[1122] = lut_1122_ff;
    end
    else begin : no_ff_1122
        assign out_data[1122] = lut_1122_out;
    end
    endgenerate
    
    
    
    // LUT : 1123
    wire [63:0] lut_1123_table = 64'b1111101110111011111110111011001110111011001100111011001100110010;
    wire [5:0] lut_1123_select = {
                             in_data[230],
                             in_data[198],
                             in_data[306],
                             in_data[219],
                             in_data[707],
                             in_data[536]};
    
    wire lut_1123_out = lut_1123_table[lut_1123_select];
    
    generate
    if ( USE_REG ) begin : ff_1123
        reg   lut_1123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1123_ff <= lut_1123_out;
            end
        end
        
        assign out_data[1123] = lut_1123_ff;
    end
    else begin : no_ff_1123
        assign out_data[1123] = lut_1123_out;
    end
    endgenerate
    
    
    
    // LUT : 1124
    wire [63:0] lut_1124_table = 64'b1111111101010101111111110111010111010101010100001111010101010001;
    wire [5:0] lut_1124_select = {
                             in_data[283],
                             in_data[471],
                             in_data[386],
                             in_data[359],
                             in_data[176],
                             in_data[215]};
    
    wire lut_1124_out = lut_1124_table[lut_1124_select];
    
    generate
    if ( USE_REG ) begin : ff_1124
        reg   lut_1124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1124_ff <= lut_1124_out;
            end
        end
        
        assign out_data[1124] = lut_1124_ff;
    end
    else begin : no_ff_1124
        assign out_data[1124] = lut_1124_out;
    end
    endgenerate
    
    
    
    // LUT : 1125
    wire [63:0] lut_1125_table = 64'b1111111111111111111111111111111111001100000000001100110000000000;
    wire [5:0] lut_1125_select = {
                             in_data[431],
                             in_data[2],
                             in_data[607],
                             in_data[562],
                             in_data[356],
                             in_data[76]};
    
    wire lut_1125_out = lut_1125_table[lut_1125_select];
    
    generate
    if ( USE_REG ) begin : ff_1125
        reg   lut_1125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1125_ff <= lut_1125_out;
            end
        end
        
        assign out_data[1125] = lut_1125_ff;
    end
    else begin : no_ff_1125
        assign out_data[1125] = lut_1125_out;
    end
    endgenerate
    
    
    
    // LUT : 1126
    wire [63:0] lut_1126_table = 64'b1111000011110000111100101111001011110011111100001111001111110011;
    wire [5:0] lut_1126_select = {
                             in_data[165],
                             in_data[409],
                             in_data[530],
                             in_data[622],
                             in_data[719],
                             in_data[583]};
    
    wire lut_1126_out = lut_1126_table[lut_1126_select];
    
    generate
    if ( USE_REG ) begin : ff_1126
        reg   lut_1126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1126_ff <= lut_1126_out;
            end
        end
        
        assign out_data[1126] = lut_1126_ff;
    end
    else begin : no_ff_1126
        assign out_data[1126] = lut_1126_out;
    end
    endgenerate
    
    
    
    // LUT : 1127
    wire [63:0] lut_1127_table = 64'b0101111101001101010111010000010000001111010111110101110101010101;
    wire [5:0] lut_1127_select = {
                             in_data[271],
                             in_data[122],
                             in_data[604],
                             in_data[211],
                             in_data[96],
                             in_data[564]};
    
    wire lut_1127_out = lut_1127_table[lut_1127_select];
    
    generate
    if ( USE_REG ) begin : ff_1127
        reg   lut_1127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1127_ff <= lut_1127_out;
            end
        end
        
        assign out_data[1127] = lut_1127_ff;
    end
    else begin : no_ff_1127
        assign out_data[1127] = lut_1127_out;
    end
    endgenerate
    
    
    
    // LUT : 1128
    wire [63:0] lut_1128_table = 64'b1111111111111111101110111111111110111011101110110010001000100010;
    wire [5:0] lut_1128_select = {
                             in_data[689],
                             in_data[276],
                             in_data[759],
                             in_data[588],
                             in_data[555],
                             in_data[255]};
    
    wire lut_1128_out = lut_1128_table[lut_1128_select];
    
    generate
    if ( USE_REG ) begin : ff_1128
        reg   lut_1128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1128_ff <= lut_1128_out;
            end
        end
        
        assign out_data[1128] = lut_1128_ff;
    end
    else begin : no_ff_1128
        assign out_data[1128] = lut_1128_out;
    end
    endgenerate
    
    
    
    // LUT : 1129
    wire [63:0] lut_1129_table = 64'b0001000000010001000001010000110100000000010101000000010100001101;
    wire [5:0] lut_1129_select = {
                             in_data[58],
                             in_data[600],
                             in_data[72],
                             in_data[377],
                             in_data[438],
                             in_data[538]};
    
    wire lut_1129_out = lut_1129_table[lut_1129_select];
    
    generate
    if ( USE_REG ) begin : ff_1129
        reg   lut_1129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1129_ff <= lut_1129_out;
            end
        end
        
        assign out_data[1129] = lut_1129_ff;
    end
    else begin : no_ff_1129
        assign out_data[1129] = lut_1129_out;
    end
    endgenerate
    
    
    
    // LUT : 1130
    wire [63:0] lut_1130_table = 64'b0000110011111111101011111111111100000000110011000000000011001110;
    wire [5:0] lut_1130_select = {
                             in_data[175],
                             in_data[748],
                             in_data[385],
                             in_data[224],
                             in_data[489],
                             in_data[23]};
    
    wire lut_1130_out = lut_1130_table[lut_1130_select];
    
    generate
    if ( USE_REG ) begin : ff_1130
        reg   lut_1130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1130_ff <= lut_1130_out;
            end
        end
        
        assign out_data[1130] = lut_1130_ff;
    end
    else begin : no_ff_1130
        assign out_data[1130] = lut_1130_out;
    end
    endgenerate
    
    
    
    // LUT : 1131
    wire [63:0] lut_1131_table = 64'b0011001000110011001100110011001111111110111111101111110011111100;
    wire [5:0] lut_1131_select = {
                             in_data[205],
                             in_data[769],
                             in_data[699],
                             in_data[526],
                             in_data[661],
                             in_data[407]};
    
    wire lut_1131_out = lut_1131_table[lut_1131_select];
    
    generate
    if ( USE_REG ) begin : ff_1131
        reg   lut_1131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1131_ff <= lut_1131_out;
            end
        end
        
        assign out_data[1131] = lut_1131_ff;
    end
    else begin : no_ff_1131
        assign out_data[1131] = lut_1131_out;
    end
    endgenerate
    
    
    
    // LUT : 1132
    wire [63:0] lut_1132_table = 64'b1011111010111000111111101111100010111110101110001111111011111000;
    wire [5:0] lut_1132_select = {
                             in_data[52],
                             in_data[14],
                             in_data[346],
                             in_data[400],
                             in_data[402],
                             in_data[677]};
    
    wire lut_1132_out = lut_1132_table[lut_1132_select];
    
    generate
    if ( USE_REG ) begin : ff_1132
        reg   lut_1132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1132_ff <= lut_1132_out;
            end
        end
        
        assign out_data[1132] = lut_1132_ff;
    end
    else begin : no_ff_1132
        assign out_data[1132] = lut_1132_out;
    end
    endgenerate
    
    
    
    // LUT : 1133
    wire [63:0] lut_1133_table = 64'b0000010001001100000001000100110000000100010011000000000001001100;
    wire [5:0] lut_1133_select = {
                             in_data[455],
                             in_data[28],
                             in_data[705],
                             in_data[423],
                             in_data[414],
                             in_data[338]};
    
    wire lut_1133_out = lut_1133_table[lut_1133_select];
    
    generate
    if ( USE_REG ) begin : ff_1133
        reg   lut_1133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1133_ff <= lut_1133_out;
            end
        end
        
        assign out_data[1133] = lut_1133_ff;
    end
    else begin : no_ff_1133
        assign out_data[1133] = lut_1133_out;
    end
    endgenerate
    
    
    
    // LUT : 1134
    wire [63:0] lut_1134_table = 64'b1111111111111111111111111111111111111111111111111111101111111010;
    wire [5:0] lut_1134_select = {
                             in_data[422],
                             in_data[254],
                             in_data[732],
                             in_data[425],
                             in_data[20],
                             in_data[117]};
    
    wire lut_1134_out = lut_1134_table[lut_1134_select];
    
    generate
    if ( USE_REG ) begin : ff_1134
        reg   lut_1134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1134_ff <= lut_1134_out;
            end
        end
        
        assign out_data[1134] = lut_1134_ff;
    end
    else begin : no_ff_1134
        assign out_data[1134] = lut_1134_out;
    end
    endgenerate
    
    
    
    // LUT : 1135
    wire [63:0] lut_1135_table = 64'b0011101100101011001111110000110000111011001110111011111100001100;
    wire [5:0] lut_1135_select = {
                             in_data[758],
                             in_data[327],
                             in_data[623],
                             in_data[174],
                             in_data[299],
                             in_data[295]};
    
    wire lut_1135_out = lut_1135_table[lut_1135_select];
    
    generate
    if ( USE_REG ) begin : ff_1135
        reg   lut_1135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1135_ff <= lut_1135_out;
            end
        end
        
        assign out_data[1135] = lut_1135_ff;
    end
    else begin : no_ff_1135
        assign out_data[1135] = lut_1135_out;
    end
    endgenerate
    
    
    
    // LUT : 1136
    wire [63:0] lut_1136_table = 64'b1100110011001100110011001100110011111111110011111111111111001110;
    wire [5:0] lut_1136_select = {
                             in_data[118],
                             in_data[503],
                             in_data[107],
                             in_data[671],
                             in_data[94],
                             in_data[17]};
    
    wire lut_1136_out = lut_1136_table[lut_1136_select];
    
    generate
    if ( USE_REG ) begin : ff_1136
        reg   lut_1136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1136_ff <= lut_1136_out;
            end
        end
        
        assign out_data[1136] = lut_1136_ff;
    end
    else begin : no_ff_1136
        assign out_data[1136] = lut_1136_out;
    end
    endgenerate
    
    
    
    // LUT : 1137
    wire [63:0] lut_1137_table = 64'b0000000000000000000010110000111111111111111111110000111100101111;
    wire [5:0] lut_1137_select = {
                             in_data[570],
                             in_data[485],
                             in_data[83],
                             in_data[602],
                             in_data[67],
                             in_data[228]};
    
    wire lut_1137_out = lut_1137_table[lut_1137_select];
    
    generate
    if ( USE_REG ) begin : ff_1137
        reg   lut_1137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1137_ff <= lut_1137_out;
            end
        end
        
        assign out_data[1137] = lut_1137_ff;
    end
    else begin : no_ff_1137
        assign out_data[1137] = lut_1137_out;
    end
    endgenerate
    
    
    
    // LUT : 1138
    wire [63:0] lut_1138_table = 64'b1111111110100000111111111010000011111111101010001111111111101000;
    wire [5:0] lut_1138_select = {
                             in_data[80],
                             in_data[724],
                             in_data[301],
                             in_data[287],
                             in_data[465],
                             in_data[618]};
    
    wire lut_1138_out = lut_1138_table[lut_1138_select];
    
    generate
    if ( USE_REG ) begin : ff_1138
        reg   lut_1138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1138_ff <= lut_1138_out;
            end
        end
        
        assign out_data[1138] = lut_1138_ff;
    end
    else begin : no_ff_1138
        assign out_data[1138] = lut_1138_out;
    end
    endgenerate
    
    
    
    // LUT : 1139
    wire [63:0] lut_1139_table = 64'b0000000010101010100010001110111000000000101010101010101011101110;
    wire [5:0] lut_1139_select = {
                             in_data[781],
                             in_data[662],
                             in_data[404],
                             in_data[447],
                             in_data[229],
                             in_data[234]};
    
    wire lut_1139_out = lut_1139_table[lut_1139_select];
    
    generate
    if ( USE_REG ) begin : ff_1139
        reg   lut_1139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1139_ff <= lut_1139_out;
            end
        end
        
        assign out_data[1139] = lut_1139_ff;
    end
    else begin : no_ff_1139
        assign out_data[1139] = lut_1139_out;
    end
    endgenerate
    
    
    
    // LUT : 1140
    wire [63:0] lut_1140_table = 64'b1111111111111111111111111111111100110111010011010001000101000100;
    wire [5:0] lut_1140_select = {
                             in_data[130],
                             in_data[173],
                             in_data[638],
                             in_data[141],
                             in_data[180],
                             in_data[360]};
    
    wire lut_1140_out = lut_1140_table[lut_1140_select];
    
    generate
    if ( USE_REG ) begin : ff_1140
        reg   lut_1140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1140_ff <= lut_1140_out;
            end
        end
        
        assign out_data[1140] = lut_1140_ff;
    end
    else begin : no_ff_1140
        assign out_data[1140] = lut_1140_out;
    end
    endgenerate
    
    
    
    // LUT : 1141
    wire [63:0] lut_1141_table = 64'b1111101011110111111010100101000011111111111111111010101011111111;
    wire [5:0] lut_1141_select = {
                             in_data[243],
                             in_data[720],
                             in_data[571],
                             in_data[341],
                             in_data[456],
                             in_data[654]};
    
    wire lut_1141_out = lut_1141_table[lut_1141_select];
    
    generate
    if ( USE_REG ) begin : ff_1141
        reg   lut_1141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1141_ff <= lut_1141_out;
            end
        end
        
        assign out_data[1141] = lut_1141_ff;
    end
    else begin : no_ff_1141
        assign out_data[1141] = lut_1141_out;
    end
    endgenerate
    
    
    
    // LUT : 1142
    wire [63:0] lut_1142_table = 64'b1111111111111111101010101010101011111111111111111111101011111011;
    wire [5:0] lut_1142_select = {
                             in_data[381],
                             in_data[461],
                             in_data[695],
                             in_data[676],
                             in_data[613],
                             in_data[120]};
    
    wire lut_1142_out = lut_1142_table[lut_1142_select];
    
    generate
    if ( USE_REG ) begin : ff_1142
        reg   lut_1142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1142_ff <= lut_1142_out;
            end
        end
        
        assign out_data[1142] = lut_1142_ff;
    end
    else begin : no_ff_1142
        assign out_data[1142] = lut_1142_out;
    end
    endgenerate
    
    
    
    // LUT : 1143
    wire [63:0] lut_1143_table = 64'b0000000000000000111111111111111100000000000000001010101011111111;
    wire [5:0] lut_1143_select = {
                             in_data[270],
                             in_data[350],
                             in_data[77],
                             in_data[5],
                             in_data[540],
                             in_data[740]};
    
    wire lut_1143_out = lut_1143_table[lut_1143_select];
    
    generate
    if ( USE_REG ) begin : ff_1143
        reg   lut_1143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1143_ff <= lut_1143_out;
            end
        end
        
        assign out_data[1143] = lut_1143_ff;
    end
    else begin : no_ff_1143
        assign out_data[1143] = lut_1143_out;
    end
    endgenerate
    
    
    
    // LUT : 1144
    wire [63:0] lut_1144_table = 64'b0000000000000000000000000000000000000000000000000000001100000011;
    wire [5:0] lut_1144_select = {
                             in_data[278],
                             in_data[253],
                             in_data[761],
                             in_data[333],
                             in_data[146],
                             in_data[110]};
    
    wire lut_1144_out = lut_1144_table[lut_1144_select];
    
    generate
    if ( USE_REG ) begin : ff_1144
        reg   lut_1144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1144_ff <= lut_1144_out;
            end
        end
        
        assign out_data[1144] = lut_1144_ff;
    end
    else begin : no_ff_1144
        assign out_data[1144] = lut_1144_out;
    end
    endgenerate
    
    
    
    // LUT : 1145
    wire [63:0] lut_1145_table = 64'b0000000000000000000100000001000011111111111111111111111111111111;
    wire [5:0] lut_1145_select = {
                             in_data[353],
                             in_data[767],
                             in_data[730],
                             in_data[612],
                             in_data[620],
                             in_data[655]};
    
    wire lut_1145_out = lut_1145_table[lut_1145_select];
    
    generate
    if ( USE_REG ) begin : ff_1145
        reg   lut_1145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1145_ff <= lut_1145_out;
            end
        end
        
        assign out_data[1145] = lut_1145_ff;
    end
    else begin : no_ff_1145
        assign out_data[1145] = lut_1145_out;
    end
    endgenerate
    
    
    
    // LUT : 1146
    wire [63:0] lut_1146_table = 64'b0101000001010000110100000101000000000000110101010100000011110101;
    wire [5:0] lut_1146_select = {
                             in_data[257],
                             in_data[196],
                             in_data[344],
                             in_data[630],
                             in_data[64],
                             in_data[249]};
    
    wire lut_1146_out = lut_1146_table[lut_1146_select];
    
    generate
    if ( USE_REG ) begin : ff_1146
        reg   lut_1146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1146_ff <= lut_1146_out;
            end
        end
        
        assign out_data[1146] = lut_1146_ff;
    end
    else begin : no_ff_1146
        assign out_data[1146] = lut_1146_out;
    end
    endgenerate
    
    
    
    // LUT : 1147
    wire [63:0] lut_1147_table = 64'b1101000100000000111101010000000011010001000000001111010100000000;
    wire [5:0] lut_1147_select = {
                             in_data[106],
                             in_data[609],
                             in_data[320],
                             in_data[332],
                             in_data[275],
                             in_data[710]};
    
    wire lut_1147_out = lut_1147_table[lut_1147_select];
    
    generate
    if ( USE_REG ) begin : ff_1147
        reg   lut_1147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1147_ff <= lut_1147_out;
            end
        end
        
        assign out_data[1147] = lut_1147_ff;
    end
    else begin : no_ff_1147
        assign out_data[1147] = lut_1147_out;
    end
    endgenerate
    
    
    
    // LUT : 1148
    wire [63:0] lut_1148_table = 64'b1111111111111111111111111111111111111111111111110000101000001110;
    wire [5:0] lut_1148_select = {
                             in_data[718],
                             in_data[649],
                             in_data[448],
                             in_data[192],
                             in_data[308],
                             in_data[682]};
    
    wire lut_1148_out = lut_1148_table[lut_1148_select];
    
    generate
    if ( USE_REG ) begin : ff_1148
        reg   lut_1148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1148_ff <= lut_1148_out;
            end
        end
        
        assign out_data[1148] = lut_1148_ff;
    end
    else begin : no_ff_1148
        assign out_data[1148] = lut_1148_out;
    end
    endgenerate
    
    
    
    // LUT : 1149
    wire [63:0] lut_1149_table = 64'b0000100011111111000010001111111100001000101011100000100010101111;
    wire [5:0] lut_1149_select = {
                             in_data[241],
                             in_data[251],
                             in_data[525],
                             in_data[221],
                             in_data[145],
                             in_data[668]};
    
    wire lut_1149_out = lut_1149_table[lut_1149_select];
    
    generate
    if ( USE_REG ) begin : ff_1149
        reg   lut_1149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1149_ff <= lut_1149_out;
            end
        end
        
        assign out_data[1149] = lut_1149_ff;
    end
    else begin : no_ff_1149
        assign out_data[1149] = lut_1149_out;
    end
    endgenerate
    
    
    
    // LUT : 1150
    wire [63:0] lut_1150_table = 64'b0101000001110000011100000111000011110000111100001111000011110000;
    wire [5:0] lut_1150_select = {
                             in_data[563],
                             in_data[171],
                             in_data[282],
                             in_data[634],
                             in_data[374],
                             in_data[766]};
    
    wire lut_1150_out = lut_1150_table[lut_1150_select];
    
    generate
    if ( USE_REG ) begin : ff_1150
        reg   lut_1150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1150_ff <= lut_1150_out;
            end
        end
        
        assign out_data[1150] = lut_1150_ff;
    end
    else begin : no_ff_1150
        assign out_data[1150] = lut_1150_out;
    end
    endgenerate
    
    
    
    // LUT : 1151
    wire [63:0] lut_1151_table = 64'b1111000011110100111100001111000011110100111101001111000011110000;
    wire [5:0] lut_1151_select = {
                             in_data[755],
                             in_data[532],
                             in_data[445],
                             in_data[544],
                             in_data[481],
                             in_data[608]};
    
    wire lut_1151_out = lut_1151_table[lut_1151_select];
    
    generate
    if ( USE_REG ) begin : ff_1151
        reg   lut_1151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1151_ff <= lut_1151_out;
            end
        end
        
        assign out_data[1151] = lut_1151_ff;
    end
    else begin : no_ff_1151
        assign out_data[1151] = lut_1151_out;
    end
    endgenerate
    
    
    
    // LUT : 1152
    wire [63:0] lut_1152_table = 64'b0101000001010100011101010111010111010000110100001111111111111111;
    wire [5:0] lut_1152_select = {
                             in_data[355],
                             in_data[491],
                             in_data[86],
                             in_data[500],
                             in_data[509],
                             in_data[665]};
    
    wire lut_1152_out = lut_1152_table[lut_1152_select];
    
    generate
    if ( USE_REG ) begin : ff_1152
        reg   lut_1152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1152_ff <= lut_1152_out;
            end
        end
        
        assign out_data[1152] = lut_1152_ff;
    end
    else begin : no_ff_1152
        assign out_data[1152] = lut_1152_out;
    end
    endgenerate
    
    
    
    // LUT : 1153
    wire [63:0] lut_1153_table = 64'b1011111110111111001100110011001100111111001111110000001100100011;
    wire [5:0] lut_1153_select = {
                             in_data[313],
                             in_data[584],
                             in_data[71],
                             in_data[220],
                             in_data[541],
                             in_data[628]};
    
    wire lut_1153_out = lut_1153_table[lut_1153_select];
    
    generate
    if ( USE_REG ) begin : ff_1153
        reg   lut_1153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1153_ff <= lut_1153_out;
            end
        end
        
        assign out_data[1153] = lut_1153_ff;
    end
    else begin : no_ff_1153
        assign out_data[1153] = lut_1153_out;
    end
    endgenerate
    
    
    
    // LUT : 1154
    wire [63:0] lut_1154_table = 64'b0000000000000000001100001111000000000000001000001111000011110000;
    wire [5:0] lut_1154_select = {
                             in_data[475],
                             in_data[302],
                             in_data[501],
                             in_data[656],
                             in_data[451],
                             in_data[672]};
    
    wire lut_1154_out = lut_1154_table[lut_1154_select];
    
    generate
    if ( USE_REG ) begin : ff_1154
        reg   lut_1154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1154_ff <= lut_1154_out;
            end
        end
        
        assign out_data[1154] = lut_1154_ff;
    end
    else begin : no_ff_1154
        assign out_data[1154] = lut_1154_out;
    end
    endgenerate
    
    
    
    // LUT : 1155
    wire [63:0] lut_1155_table = 64'b0000000000001111000000000000111100000010000000000000001000000000;
    wire [5:0] lut_1155_select = {
                             in_data[406],
                             in_data[51],
                             in_data[412],
                             in_data[305],
                             in_data[472],
                             in_data[151]};
    
    wire lut_1155_out = lut_1155_table[lut_1155_select];
    
    generate
    if ( USE_REG ) begin : ff_1155
        reg   lut_1155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1155_ff <= lut_1155_out;
            end
        end
        
        assign out_data[1155] = lut_1155_ff;
    end
    else begin : no_ff_1155
        assign out_data[1155] = lut_1155_out;
    end
    endgenerate
    
    
    
    // LUT : 1156
    wire [63:0] lut_1156_table = 64'b1111111111111111110111011101111111011101110111010100010001000100;
    wire [5:0] lut_1156_select = {
                             in_data[637],
                             in_data[119],
                             in_data[777],
                             in_data[79],
                             in_data[370],
                             in_data[136]};
    
    wire lut_1156_out = lut_1156_table[lut_1156_select];
    
    generate
    if ( USE_REG ) begin : ff_1156
        reg   lut_1156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1156_ff <= lut_1156_out;
            end
        end
        
        assign out_data[1156] = lut_1156_ff;
    end
    else begin : no_ff_1156
        assign out_data[1156] = lut_1156_out;
    end
    endgenerate
    
    
    
    // LUT : 1157
    wire [63:0] lut_1157_table = 64'b1111111111111111111111111111111111111111111111111111111111111010;
    wire [5:0] lut_1157_select = {
                             in_data[193],
                             in_data[75],
                             in_data[103],
                             in_data[191],
                             in_data[701],
                             in_data[125]};
    
    wire lut_1157_out = lut_1157_table[lut_1157_select];
    
    generate
    if ( USE_REG ) begin : ff_1157
        reg   lut_1157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1157_ff <= lut_1157_out;
            end
        end
        
        assign out_data[1157] = lut_1157_ff;
    end
    else begin : no_ff_1157
        assign out_data[1157] = lut_1157_out;
    end
    endgenerate
    
    
    
    // LUT : 1158
    wire [63:0] lut_1158_table = 64'b1101111111001111110011110100111111000000111111110000000011111111;
    wire [5:0] lut_1158_select = {
                             in_data[272],
                             in_data[142],
                             in_data[267],
                             in_data[454],
                             in_data[389],
                             in_data[586]};
    
    wire lut_1158_out = lut_1158_table[lut_1158_select];
    
    generate
    if ( USE_REG ) begin : ff_1158
        reg   lut_1158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1158_ff <= lut_1158_out;
            end
        end
        
        assign out_data[1158] = lut_1158_ff;
    end
    else begin : no_ff_1158
        assign out_data[1158] = lut_1158_out;
    end
    endgenerate
    
    
    
    // LUT : 1159
    wire [63:0] lut_1159_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1159_select = {
                             in_data[337],
                             in_data[7],
                             in_data[108],
                             in_data[578],
                             in_data[231],
                             in_data[617]};
    
    wire lut_1159_out = lut_1159_table[lut_1159_select];
    
    generate
    if ( USE_REG ) begin : ff_1159
        reg   lut_1159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1159_ff <= lut_1159_out;
            end
        end
        
        assign out_data[1159] = lut_1159_ff;
    end
    else begin : no_ff_1159
        assign out_data[1159] = lut_1159_out;
    end
    endgenerate
    
    
    
    // LUT : 1160
    wire [63:0] lut_1160_table = 64'b0000000000000000000000000000111100000000000000000000000000001111;
    wire [5:0] lut_1160_select = {
                             in_data[18],
                             in_data[194],
                             in_data[102],
                             in_data[747],
                             in_data[365],
                             in_data[195]};
    
    wire lut_1160_out = lut_1160_table[lut_1160_select];
    
    generate
    if ( USE_REG ) begin : ff_1160
        reg   lut_1160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1160_ff <= lut_1160_out;
            end
        end
        
        assign out_data[1160] = lut_1160_ff;
    end
    else begin : no_ff_1160
        assign out_data[1160] = lut_1160_out;
    end
    endgenerate
    
    
    
    // LUT : 1161
    wire [63:0] lut_1161_table = 64'b0010001100100011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1161_select = {
                             in_data[577],
                             in_data[366],
                             in_data[647],
                             in_data[560],
                             in_data[624],
                             in_data[66]};
    
    wire lut_1161_out = lut_1161_table[lut_1161_select];
    
    generate
    if ( USE_REG ) begin : ff_1161
        reg   lut_1161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1161_ff <= lut_1161_out;
            end
        end
        
        assign out_data[1161] = lut_1161_ff;
    end
    else begin : no_ff_1161
        assign out_data[1161] = lut_1161_out;
    end
    endgenerate
    
    
    
    // LUT : 1162
    wire [63:0] lut_1162_table = 64'b0000000000000000000000000000000000000001000000010000000100000001;
    wire [5:0] lut_1162_select = {
                             in_data[746],
                             in_data[53],
                             in_data[450],
                             in_data[129],
                             in_data[124],
                             in_data[683]};
    
    wire lut_1162_out = lut_1162_table[lut_1162_select];
    
    generate
    if ( USE_REG ) begin : ff_1162
        reg   lut_1162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1162_ff <= lut_1162_out;
            end
        end
        
        assign out_data[1162] = lut_1162_ff;
    end
    else begin : no_ff_1162
        assign out_data[1162] = lut_1162_out;
    end
    endgenerate
    
    
    
    // LUT : 1163
    wire [63:0] lut_1163_table = 64'b0000101000001010000010100000101000001010101011111010101011111111;
    wire [5:0] lut_1163_select = {
                             in_data[492],
                             in_data[750],
                             in_data[296],
                             in_data[172],
                             in_data[420],
                             in_data[330]};
    
    wire lut_1163_out = lut_1163_table[lut_1163_select];
    
    generate
    if ( USE_REG ) begin : ff_1163
        reg   lut_1163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1163_ff <= lut_1163_out;
            end
        end
        
        assign out_data[1163] = lut_1163_ff;
    end
    else begin : no_ff_1163
        assign out_data[1163] = lut_1163_out;
    end
    endgenerate
    
    
    
    // LUT : 1164
    wire [63:0] lut_1164_table = 64'b0101010101010101000000000101010001010101010101010000000000000000;
    wire [5:0] lut_1164_select = {
                             in_data[522],
                             in_data[575],
                             in_data[743],
                             in_data[55],
                             in_data[782],
                             in_data[687]};
    
    wire lut_1164_out = lut_1164_table[lut_1164_select];
    
    generate
    if ( USE_REG ) begin : ff_1164
        reg   lut_1164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1164_ff <= lut_1164_out;
            end
        end
        
        assign out_data[1164] = lut_1164_ff;
    end
    else begin : no_ff_1164
        assign out_data[1164] = lut_1164_out;
    end
    endgenerate
    
    
    
    // LUT : 1165
    wire [63:0] lut_1165_table = 64'b1010000010101010101000101010101001010000111101000101000011110100;
    wire [5:0] lut_1165_select = {
                             in_data[553],
                             in_data[3],
                             in_data[199],
                             in_data[499],
                             in_data[185],
                             in_data[517]};
    
    wire lut_1165_out = lut_1165_table[lut_1165_select];
    
    generate
    if ( USE_REG ) begin : ff_1165
        reg   lut_1165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1165_ff <= lut_1165_out;
            end
        end
        
        assign out_data[1165] = lut_1165_ff;
    end
    else begin : no_ff_1165
        assign out_data[1165] = lut_1165_out;
    end
    endgenerate
    
    
    
    // LUT : 1166
    wire [63:0] lut_1166_table = 64'b1111111111111111111111111111111111111111101110111111111110111011;
    wire [5:0] lut_1166_select = {
                             in_data[619],
                             in_data[42],
                             in_data[90],
                             in_data[4],
                             in_data[539],
                             in_data[69]};
    
    wire lut_1166_out = lut_1166_table[lut_1166_select];
    
    generate
    if ( USE_REG ) begin : ff_1166
        reg   lut_1166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1166_ff <= lut_1166_out;
            end
        end
        
        assign out_data[1166] = lut_1166_ff;
    end
    else begin : no_ff_1166
        assign out_data[1166] = lut_1166_out;
    end
    endgenerate
    
    
    
    // LUT : 1167
    wire [63:0] lut_1167_table = 64'b1111000010110000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1167_select = {
                             in_data[403],
                             in_data[242],
                             in_data[335],
                             in_data[735],
                             in_data[533],
                             in_data[39]};
    
    wire lut_1167_out = lut_1167_table[lut_1167_select];
    
    generate
    if ( USE_REG ) begin : ff_1167
        reg   lut_1167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1167_ff <= lut_1167_out;
            end
        end
        
        assign out_data[1167] = lut_1167_ff;
    end
    else begin : no_ff_1167
        assign out_data[1167] = lut_1167_out;
    end
    endgenerate
    
    
    
    // LUT : 1168
    wire [63:0] lut_1168_table = 64'b0000000000000101000000010000011100000000000000010000000000000001;
    wire [5:0] lut_1168_select = {
                             in_data[446],
                             in_data[168],
                             in_data[311],
                             in_data[397],
                             in_data[307],
                             in_data[742]};
    
    wire lut_1168_out = lut_1168_table[lut_1168_select];
    
    generate
    if ( USE_REG ) begin : ff_1168
        reg   lut_1168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1168_ff <= lut_1168_out;
            end
        end
        
        assign out_data[1168] = lut_1168_ff;
    end
    else begin : no_ff_1168
        assign out_data[1168] = lut_1168_out;
    end
    endgenerate
    
    
    
    // LUT : 1169
    wire [63:0] lut_1169_table = 64'b0000111100001111111111110010111100001000000000000010101000000000;
    wire [5:0] lut_1169_select = {
                             in_data[317],
                             in_data[258],
                             in_data[186],
                             in_data[162],
                             in_data[733],
                             in_data[675]};
    
    wire lut_1169_out = lut_1169_table[lut_1169_select];
    
    generate
    if ( USE_REG ) begin : ff_1169
        reg   lut_1169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1169_ff <= lut_1169_out;
            end
        end
        
        assign out_data[1169] = lut_1169_ff;
    end
    else begin : no_ff_1169
        assign out_data[1169] = lut_1169_out;
    end
    endgenerate
    
    
    
    // LUT : 1170
    wire [63:0] lut_1170_table = 64'b0011001100000000001100110000000000110011000000000011001100000000;
    wire [5:0] lut_1170_select = {
                             in_data[174],
                             in_data[69],
                             in_data[259],
                             in_data[134],
                             in_data[554],
                             in_data[115]};
    
    wire lut_1170_out = lut_1170_table[lut_1170_select];
    
    generate
    if ( USE_REG ) begin : ff_1170
        reg   lut_1170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1170_ff <= lut_1170_out;
            end
        end
        
        assign out_data[1170] = lut_1170_ff;
    end
    else begin : no_ff_1170
        assign out_data[1170] = lut_1170_out;
    end
    endgenerate
    
    
    
    // LUT : 1171
    wire [63:0] lut_1171_table = 64'b1111111111111010111111111111101011111111111110101111111111111010;
    wire [5:0] lut_1171_select = {
                             in_data[196],
                             in_data[309],
                             in_data[491],
                             in_data[423],
                             in_data[197],
                             in_data[692]};
    
    wire lut_1171_out = lut_1171_table[lut_1171_select];
    
    generate
    if ( USE_REG ) begin : ff_1171
        reg   lut_1171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1171_ff <= lut_1171_out;
            end
        end
        
        assign out_data[1171] = lut_1171_ff;
    end
    else begin : no_ff_1171
        assign out_data[1171] = lut_1171_out;
    end
    endgenerate
    
    
    
    // LUT : 1172
    wire [63:0] lut_1172_table = 64'b1111111111111100111111111111111011110011111100001111001111110000;
    wire [5:0] lut_1172_select = {
                             in_data[273],
                             in_data[114],
                             in_data[355],
                             in_data[655],
                             in_data[401],
                             in_data[704]};
    
    wire lut_1172_out = lut_1172_table[lut_1172_select];
    
    generate
    if ( USE_REG ) begin : ff_1172
        reg   lut_1172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1172_ff <= lut_1172_out;
            end
        end
        
        assign out_data[1172] = lut_1172_ff;
    end
    else begin : no_ff_1172
        assign out_data[1172] = lut_1172_out;
    end
    endgenerate
    
    
    
    // LUT : 1173
    wire [63:0] lut_1173_table = 64'b0000000000000000000000000000000000000000000100010000000000110011;
    wire [5:0] lut_1173_select = {
                             in_data[743],
                             in_data[565],
                             in_data[695],
                             in_data[139],
                             in_data[240],
                             in_data[391]};
    
    wire lut_1173_out = lut_1173_table[lut_1173_select];
    
    generate
    if ( USE_REG ) begin : ff_1173
        reg   lut_1173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1173_ff <= lut_1173_out;
            end
        end
        
        assign out_data[1173] = lut_1173_ff;
    end
    else begin : no_ff_1173
        assign out_data[1173] = lut_1173_out;
    end
    endgenerate
    
    
    
    // LUT : 1174
    wire [63:0] lut_1174_table = 64'b0000000000000000000000000000000000000000000000000010101010101011;
    wire [5:0] lut_1174_select = {
                             in_data[248],
                             in_data[742],
                             in_data[589],
                             in_data[586],
                             in_data[668],
                             in_data[389]};
    
    wire lut_1174_out = lut_1174_table[lut_1174_select];
    
    generate
    if ( USE_REG ) begin : ff_1174
        reg   lut_1174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1174_ff <= lut_1174_out;
            end
        end
        
        assign out_data[1174] = lut_1174_ff;
    end
    else begin : no_ff_1174
        assign out_data[1174] = lut_1174_out;
    end
    endgenerate
    
    
    
    // LUT : 1175
    wire [63:0] lut_1175_table = 64'b0000111100000000000011110000000000001111000000000000111100000000;
    wire [5:0] lut_1175_select = {
                             in_data[62],
                             in_data[27],
                             in_data[266],
                             in_data[592],
                             in_data[736],
                             in_data[562]};
    
    wire lut_1175_out = lut_1175_table[lut_1175_select];
    
    generate
    if ( USE_REG ) begin : ff_1175
        reg   lut_1175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1175_ff <= lut_1175_out;
            end
        end
        
        assign out_data[1175] = lut_1175_ff;
    end
    else begin : no_ff_1175
        assign out_data[1175] = lut_1175_out;
    end
    endgenerate
    
    
    
    // LUT : 1176
    wire [63:0] lut_1176_table = 64'b1111111111111111111100001111000011010101110101010000000000000000;
    wire [5:0] lut_1176_select = {
                             in_data[373],
                             in_data[241],
                             in_data[171],
                             in_data[520],
                             in_data[691],
                             in_data[576]};
    
    wire lut_1176_out = lut_1176_table[lut_1176_select];
    
    generate
    if ( USE_REG ) begin : ff_1176
        reg   lut_1176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1176_ff <= lut_1176_out;
            end
        end
        
        assign out_data[1176] = lut_1176_ff;
    end
    else begin : no_ff_1176
        assign out_data[1176] = lut_1176_out;
    end
    endgenerate
    
    
    
    // LUT : 1177
    wire [63:0] lut_1177_table = 64'b1111111100001111100011110000100011111111111111110000111000000000;
    wire [5:0] lut_1177_select = {
                             in_data[357],
                             in_data[263],
                             in_data[610],
                             in_data[416],
                             in_data[766],
                             in_data[584]};
    
    wire lut_1177_out = lut_1177_table[lut_1177_select];
    
    generate
    if ( USE_REG ) begin : ff_1177
        reg   lut_1177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1177_ff <= lut_1177_out;
            end
        end
        
        assign out_data[1177] = lut_1177_ff;
    end
    else begin : no_ff_1177
        assign out_data[1177] = lut_1177_out;
    end
    endgenerate
    
    
    
    // LUT : 1178
    wire [63:0] lut_1178_table = 64'b1111111111111111111111111111011111110101010100011111010111010000;
    wire [5:0] lut_1178_select = {
                             in_data[713],
                             in_data[694],
                             in_data[712],
                             in_data[471],
                             in_data[512],
                             in_data[333]};
    
    wire lut_1178_out = lut_1178_table[lut_1178_select];
    
    generate
    if ( USE_REG ) begin : ff_1178
        reg   lut_1178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1178_ff <= lut_1178_out;
            end
        end
        
        assign out_data[1178] = lut_1178_ff;
    end
    else begin : no_ff_1178
        assign out_data[1178] = lut_1178_out;
    end
    endgenerate
    
    
    
    // LUT : 1179
    wire [63:0] lut_1179_table = 64'b0000000000010101000001010000010100000000000001010000010101000101;
    wire [5:0] lut_1179_select = {
                             in_data[353],
                             in_data[368],
                             in_data[385],
                             in_data[414],
                             in_data[81],
                             in_data[219]};
    
    wire lut_1179_out = lut_1179_table[lut_1179_select];
    
    generate
    if ( USE_REG ) begin : ff_1179
        reg   lut_1179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1179_ff <= lut_1179_out;
            end
        end
        
        assign out_data[1179] = lut_1179_ff;
    end
    else begin : no_ff_1179
        assign out_data[1179] = lut_1179_out;
    end
    endgenerate
    
    
    
    // LUT : 1180
    wire [63:0] lut_1180_table = 64'b0000000000000000000000001100110011111110111111111111111111111111;
    wire [5:0] lut_1180_select = {
                             in_data[384],
                             in_data[518],
                             in_data[651],
                             in_data[366],
                             in_data[189],
                             in_data[530]};
    
    wire lut_1180_out = lut_1180_table[lut_1180_select];
    
    generate
    if ( USE_REG ) begin : ff_1180
        reg   lut_1180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1180_ff <= lut_1180_out;
            end
        end
        
        assign out_data[1180] = lut_1180_ff;
    end
    else begin : no_ff_1180
        assign out_data[1180] = lut_1180_out;
    end
    endgenerate
    
    
    
    // LUT : 1181
    wire [63:0] lut_1181_table = 64'b0000000000000000000000000000000000000011000000110000001000000001;
    wire [5:0] lut_1181_select = {
                             in_data[583],
                             in_data[761],
                             in_data[33],
                             in_data[479],
                             in_data[776],
                             in_data[560]};
    
    wire lut_1181_out = lut_1181_table[lut_1181_select];
    
    generate
    if ( USE_REG ) begin : ff_1181
        reg   lut_1181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1181_ff <= lut_1181_out;
            end
        end
        
        assign out_data[1181] = lut_1181_ff;
    end
    else begin : no_ff_1181
        assign out_data[1181] = lut_1181_out;
    end
    endgenerate
    
    
    
    // LUT : 1182
    wire [63:0] lut_1182_table = 64'b0000000000000001000100010001000100000000000001000100110101011101;
    wire [5:0] lut_1182_select = {
                             in_data[186],
                             in_data[539],
                             in_data[758],
                             in_data[67],
                             in_data[632],
                             in_data[468]};
    
    wire lut_1182_out = lut_1182_table[lut_1182_select];
    
    generate
    if ( USE_REG ) begin : ff_1182
        reg   lut_1182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1182_ff <= lut_1182_out;
            end
        end
        
        assign out_data[1182] = lut_1182_ff;
    end
    else begin : no_ff_1182
        assign out_data[1182] = lut_1182_out;
    end
    endgenerate
    
    
    
    // LUT : 1183
    wire [63:0] lut_1183_table = 64'b1100000011111101111100001111110001000000111111000100000011111100;
    wire [5:0] lut_1183_select = {
                             in_data[77],
                             in_data[505],
                             in_data[262],
                             in_data[571],
                             in_data[101],
                             in_data[675]};
    
    wire lut_1183_out = lut_1183_table[lut_1183_select];
    
    generate
    if ( USE_REG ) begin : ff_1183
        reg   lut_1183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1183_ff <= lut_1183_out;
            end
        end
        
        assign out_data[1183] = lut_1183_ff;
    end
    else begin : no_ff_1183
        assign out_data[1183] = lut_1183_out;
    end
    endgenerate
    
    
    
    // LUT : 1184
    wire [63:0] lut_1184_table = 64'b1111111111111111111100001111000011111111111111111111000011111000;
    wire [5:0] lut_1184_select = {
                             in_data[84],
                             in_data[715],
                             in_data[528],
                             in_data[621],
                             in_data[328],
                             in_data[32]};
    
    wire lut_1184_out = lut_1184_table[lut_1184_select];
    
    generate
    if ( USE_REG ) begin : ff_1184
        reg   lut_1184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1184_ff <= lut_1184_out;
            end
        end
        
        assign out_data[1184] = lut_1184_ff;
    end
    else begin : no_ff_1184
        assign out_data[1184] = lut_1184_out;
    end
    endgenerate
    
    
    
    // LUT : 1185
    wire [63:0] lut_1185_table = 64'b1111111100000000000000000000000000100011111111110000000010111011;
    wire [5:0] lut_1185_select = {
                             in_data[511],
                             in_data[236],
                             in_data[456],
                             in_data[723],
                             in_data[753],
                             in_data[40]};
    
    wire lut_1185_out = lut_1185_table[lut_1185_select];
    
    generate
    if ( USE_REG ) begin : ff_1185
        reg   lut_1185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1185_ff <= lut_1185_out;
            end
        end
        
        assign out_data[1185] = lut_1185_ff;
    end
    else begin : no_ff_1185
        assign out_data[1185] = lut_1185_out;
    end
    endgenerate
    
    
    
    // LUT : 1186
    wire [63:0] lut_1186_table = 64'b0000000000000000110111011000100000000000000000001101110110001001;
    wire [5:0] lut_1186_select = {
                             in_data[644],
                             in_data[102],
                             in_data[212],
                             in_data[167],
                             in_data[161],
                             in_data[525]};
    
    wire lut_1186_out = lut_1186_table[lut_1186_select];
    
    generate
    if ( USE_REG ) begin : ff_1186
        reg   lut_1186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1186_ff <= lut_1186_out;
            end
        end
        
        assign out_data[1186] = lut_1186_ff;
    end
    else begin : no_ff_1186
        assign out_data[1186] = lut_1186_out;
    end
    endgenerate
    
    
    
    // LUT : 1187
    wire [63:0] lut_1187_table = 64'b0000000011101000001100001111110000000000111011000011000011111110;
    wire [5:0] lut_1187_select = {
                             in_data[645],
                             in_data[75],
                             in_data[648],
                             in_data[748],
                             in_data[654],
                             in_data[250]};
    
    wire lut_1187_out = lut_1187_table[lut_1187_select];
    
    generate
    if ( USE_REG ) begin : ff_1187
        reg   lut_1187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1187_ff <= lut_1187_out;
            end
        end
        
        assign out_data[1187] = lut_1187_ff;
    end
    else begin : no_ff_1187
        assign out_data[1187] = lut_1187_out;
    end
    endgenerate
    
    
    
    // LUT : 1188
    wire [63:0] lut_1188_table = 64'b0011111100000000101111110000000011111111000000001111111100110000;
    wire [5:0] lut_1188_select = {
                             in_data[163],
                             in_data[740],
                             in_data[329],
                             in_data[153],
                             in_data[182],
                             in_data[697]};
    
    wire lut_1188_out = lut_1188_table[lut_1188_select];
    
    generate
    if ( USE_REG ) begin : ff_1188
        reg   lut_1188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1188_ff <= lut_1188_out;
            end
        end
        
        assign out_data[1188] = lut_1188_ff;
    end
    else begin : no_ff_1188
        assign out_data[1188] = lut_1188_out;
    end
    endgenerate
    
    
    
    // LUT : 1189
    wire [63:0] lut_1189_table = 64'b0101010101010101111111111111111100000000000000000000000000000000;
    wire [5:0] lut_1189_select = {
                             in_data[687],
                             in_data[650],
                             in_data[59],
                             in_data[726],
                             in_data[278],
                             in_data[507]};
    
    wire lut_1189_out = lut_1189_table[lut_1189_select];
    
    generate
    if ( USE_REG ) begin : ff_1189
        reg   lut_1189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1189_ff <= lut_1189_out;
            end
        end
        
        assign out_data[1189] = lut_1189_ff;
    end
    else begin : no_ff_1189
        assign out_data[1189] = lut_1189_out;
    end
    endgenerate
    
    
    
    // LUT : 1190
    wire [63:0] lut_1190_table = 64'b1111111100000000111111110101000011111111000000001111111111010000;
    wire [5:0] lut_1190_select = {
                             in_data[365],
                             in_data[46],
                             in_data[558],
                             in_data[166],
                             in_data[2],
                             in_data[419]};
    
    wire lut_1190_out = lut_1190_table[lut_1190_select];
    
    generate
    if ( USE_REG ) begin : ff_1190
        reg   lut_1190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1190_ff <= lut_1190_out;
            end
        end
        
        assign out_data[1190] = lut_1190_ff;
    end
    else begin : no_ff_1190
        assign out_data[1190] = lut_1190_out;
    end
    endgenerate
    
    
    
    // LUT : 1191
    wire [63:0] lut_1191_table = 64'b0000000101010101000001010101010100000000000101010000000000000000;
    wire [5:0] lut_1191_select = {
                             in_data[242],
                             in_data[612],
                             in_data[323],
                             in_data[253],
                             in_data[752],
                             in_data[125]};
    
    wire lut_1191_out = lut_1191_table[lut_1191_select];
    
    generate
    if ( USE_REG ) begin : ff_1191
        reg   lut_1191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1191_ff <= lut_1191_out;
            end
        end
        
        assign out_data[1191] = lut_1191_ff;
    end
    else begin : no_ff_1191
        assign out_data[1191] = lut_1191_out;
    end
    endgenerate
    
    
    
    // LUT : 1192
    wire [63:0] lut_1192_table = 64'b1010000000000000000000000000000011111000111100001111100011110000;
    wire [5:0] lut_1192_select = {
                             in_data[593],
                             in_data[763],
                             in_data[354],
                             in_data[486],
                             in_data[396],
                             in_data[737]};
    
    wire lut_1192_out = lut_1192_table[lut_1192_select];
    
    generate
    if ( USE_REG ) begin : ff_1192
        reg   lut_1192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1192_ff <= lut_1192_out;
            end
        end
        
        assign out_data[1192] = lut_1192_ff;
    end
    else begin : no_ff_1192
        assign out_data[1192] = lut_1192_out;
    end
    endgenerate
    
    
    
    // LUT : 1193
    wire [63:0] lut_1193_table = 64'b1000100010001000110110011101110110001000100010001101100011011000;
    wire [5:0] lut_1193_select = {
                             in_data[314],
                             in_data[611],
                             in_data[727],
                             in_data[113],
                             in_data[374],
                             in_data[521]};
    
    wire lut_1193_out = lut_1193_table[lut_1193_select];
    
    generate
    if ( USE_REG ) begin : ff_1193
        reg   lut_1193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1193_ff <= lut_1193_out;
            end
        end
        
        assign out_data[1193] = lut_1193_ff;
    end
    else begin : no_ff_1193
        assign out_data[1193] = lut_1193_out;
    end
    endgenerate
    
    
    
    // LUT : 1194
    wire [63:0] lut_1194_table = 64'b0000000000000000001000001111000100000000000000001010000011110101;
    wire [5:0] lut_1194_select = {
                             in_data[38],
                             in_data[538],
                             in_data[599],
                             in_data[457],
                             in_data[108],
                             in_data[487]};
    
    wire lut_1194_out = lut_1194_table[lut_1194_select];
    
    generate
    if ( USE_REG ) begin : ff_1194
        reg   lut_1194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1194_ff <= lut_1194_out;
            end
        end
        
        assign out_data[1194] = lut_1194_ff;
    end
    else begin : no_ff_1194
        assign out_data[1194] = lut_1194_out;
    end
    endgenerate
    
    
    
    // LUT : 1195
    wire [63:0] lut_1195_table = 64'b1111111111111111000000000000000010111111101111110000000000000000;
    wire [5:0] lut_1195_select = {
                             in_data[229],
                             in_data[372],
                             in_data[722],
                             in_data[405],
                             in_data[734],
                             in_data[261]};
    
    wire lut_1195_out = lut_1195_table[lut_1195_select];
    
    generate
    if ( USE_REG ) begin : ff_1195
        reg   lut_1195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1195_ff <= lut_1195_out;
            end
        end
        
        assign out_data[1195] = lut_1195_ff;
    end
    else begin : no_ff_1195
        assign out_data[1195] = lut_1195_out;
    end
    endgenerate
    
    
    
    // LUT : 1196
    wire [63:0] lut_1196_table = 64'b1101110111011111110111111111111100000100000001000100010100000101;
    wire [5:0] lut_1196_select = {
                             in_data[634],
                             in_data[567],
                             in_data[68],
                             in_data[582],
                             in_data[177],
                             in_data[294]};
    
    wire lut_1196_out = lut_1196_table[lut_1196_select];
    
    generate
    if ( USE_REG ) begin : ff_1196
        reg   lut_1196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1196_ff <= lut_1196_out;
            end
        end
        
        assign out_data[1196] = lut_1196_ff;
    end
    else begin : no_ff_1196
        assign out_data[1196] = lut_1196_out;
    end
    endgenerate
    
    
    
    // LUT : 1197
    wire [63:0] lut_1197_table = 64'b1111111111111111101111111111111110111011001100000010101000000000;
    wire [5:0] lut_1197_select = {
                             in_data[207],
                             in_data[100],
                             in_data[628],
                             in_data[246],
                             in_data[200],
                             in_data[609]};
    
    wire lut_1197_out = lut_1197_table[lut_1197_select];
    
    generate
    if ( USE_REG ) begin : ff_1197
        reg   lut_1197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1197_ff <= lut_1197_out;
            end
        end
        
        assign out_data[1197] = lut_1197_ff;
    end
    else begin : no_ff_1197
        assign out_data[1197] = lut_1197_out;
    end
    endgenerate
    
    
    
    // LUT : 1198
    wire [63:0] lut_1198_table = 64'b0000000000000000000000000000000000000101000001010000010100000101;
    wire [5:0] lut_1198_select = {
                             in_data[301],
                             in_data[307],
                             in_data[55],
                             in_data[711],
                             in_data[674],
                             in_data[346]};
    
    wire lut_1198_out = lut_1198_table[lut_1198_select];
    
    generate
    if ( USE_REG ) begin : ff_1198
        reg   lut_1198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1198_ff <= lut_1198_out;
            end
        end
        
        assign out_data[1198] = lut_1198_ff;
    end
    else begin : no_ff_1198
        assign out_data[1198] = lut_1198_out;
    end
    endgenerate
    
    
    
    // LUT : 1199
    wire [63:0] lut_1199_table = 64'b0000000000000000111100001111000001110000001100001111000011110001;
    wire [5:0] lut_1199_select = {
                             in_data[303],
                             in_data[424],
                             in_data[733],
                             in_data[536],
                             in_data[719],
                             in_data[671]};
    
    wire lut_1199_out = lut_1199_table[lut_1199_select];
    
    generate
    if ( USE_REG ) begin : ff_1199
        reg   lut_1199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1199_ff <= lut_1199_out;
            end
        end
        
        assign out_data[1199] = lut_1199_ff;
    end
    else begin : no_ff_1199
        assign out_data[1199] = lut_1199_out;
    end
    endgenerate
    
    
    
    // LUT : 1200
    wire [63:0] lut_1200_table = 64'b1111111111111111010011000100111011111111111111111100010001001000;
    wire [5:0] lut_1200_select = {
                             in_data[98],
                             in_data[325],
                             in_data[639],
                             in_data[231],
                             in_data[378],
                             in_data[496]};
    
    wire lut_1200_out = lut_1200_table[lut_1200_select];
    
    generate
    if ( USE_REG ) begin : ff_1200
        reg   lut_1200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1200_ff <= lut_1200_out;
            end
        end
        
        assign out_data[1200] = lut_1200_ff;
    end
    else begin : no_ff_1200
        assign out_data[1200] = lut_1200_out;
    end
    endgenerate
    
    
    
    // LUT : 1201
    wire [63:0] lut_1201_table = 64'b0111011101010111011101110111011100010001000100010001000100010001;
    wire [5:0] lut_1201_select = {
                             in_data[570],
                             in_data[680],
                             in_data[17],
                             in_data[308],
                             in_data[238],
                             in_data[287]};
    
    wire lut_1201_out = lut_1201_table[lut_1201_select];
    
    generate
    if ( USE_REG ) begin : ff_1201
        reg   lut_1201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1201_ff <= lut_1201_out;
            end
        end
        
        assign out_data[1201] = lut_1201_ff;
    end
    else begin : no_ff_1201
        assign out_data[1201] = lut_1201_out;
    end
    endgenerate
    
    
    
    // LUT : 1202
    wire [63:0] lut_1202_table = 64'b0000000000000000000000000000000011001100000000001100110011001100;
    wire [5:0] lut_1202_select = {
                             in_data[707],
                             in_data[202],
                             in_data[286],
                             in_data[49],
                             in_data[455],
                             in_data[58]};
    
    wire lut_1202_out = lut_1202_table[lut_1202_select];
    
    generate
    if ( USE_REG ) begin : ff_1202
        reg   lut_1202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1202_ff <= lut_1202_out;
            end
        end
        
        assign out_data[1202] = lut_1202_ff;
    end
    else begin : no_ff_1202
        assign out_data[1202] = lut_1202_out;
    end
    endgenerate
    
    
    
    // LUT : 1203
    wire [63:0] lut_1203_table = 64'b1111111111111111111110001111110011111111111111111111000011110000;
    wire [5:0] lut_1203_select = {
                             in_data[429],
                             in_data[342],
                             in_data[703],
                             in_data[320],
                             in_data[191],
                             in_data[458]};
    
    wire lut_1203_out = lut_1203_table[lut_1203_select];
    
    generate
    if ( USE_REG ) begin : ff_1203
        reg   lut_1203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1203_ff <= lut_1203_out;
            end
        end
        
        assign out_data[1203] = lut_1203_ff;
    end
    else begin : no_ff_1203
        assign out_data[1203] = lut_1203_out;
    end
    endgenerate
    
    
    
    // LUT : 1204
    wire [63:0] lut_1204_table = 64'b1111010111110000111101011111010111110101111101011111010111110001;
    wire [5:0] lut_1204_select = {
                             in_data[90],
                             in_data[201],
                             in_data[260],
                             in_data[620],
                             in_data[614],
                             in_data[497]};
    
    wire lut_1204_out = lut_1204_table[lut_1204_select];
    
    generate
    if ( USE_REG ) begin : ff_1204
        reg   lut_1204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1204_ff <= lut_1204_out;
            end
        end
        
        assign out_data[1204] = lut_1204_ff;
    end
    else begin : no_ff_1204
        assign out_data[1204] = lut_1204_out;
    end
    endgenerate
    
    
    
    // LUT : 1205
    wire [63:0] lut_1205_table = 64'b1111111101011101111111110101110111111111101010101110111010101010;
    wire [5:0] lut_1205_select = {
                             in_data[498],
                             in_data[142],
                             in_data[481],
                             in_data[701],
                             in_data[107],
                             in_data[467]};
    
    wire lut_1205_out = lut_1205_table[lut_1205_select];
    
    generate
    if ( USE_REG ) begin : ff_1205
        reg   lut_1205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1205_ff <= lut_1205_out;
            end
        end
        
        assign out_data[1205] = lut_1205_ff;
    end
    else begin : no_ff_1205
        assign out_data[1205] = lut_1205_out;
    end
    endgenerate
    
    
    
    // LUT : 1206
    wire [63:0] lut_1206_table = 64'b0000000000000000001100010011001100000000000000000011000100110011;
    wire [5:0] lut_1206_select = {
                             in_data[3],
                             in_data[176],
                             in_data[324],
                             in_data[717],
                             in_data[232],
                             in_data[624]};
    
    wire lut_1206_out = lut_1206_table[lut_1206_select];
    
    generate
    if ( USE_REG ) begin : ff_1206
        reg   lut_1206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1206_ff <= lut_1206_out;
            end
        end
        
        assign out_data[1206] = lut_1206_ff;
    end
    else begin : no_ff_1206
        assign out_data[1206] = lut_1206_out;
    end
    endgenerate
    
    
    
    // LUT : 1207
    wire [63:0] lut_1207_table = 64'b1111111111111111000000000000000010111111111111110000000000000000;
    wire [5:0] lut_1207_select = {
                             in_data[319],
                             in_data[434],
                             in_data[569],
                             in_data[223],
                             in_data[749],
                             in_data[382]};
    
    wire lut_1207_out = lut_1207_table[lut_1207_select];
    
    generate
    if ( USE_REG ) begin : ff_1207
        reg   lut_1207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1207_ff <= lut_1207_out;
            end
        end
        
        assign out_data[1207] = lut_1207_ff;
    end
    else begin : no_ff_1207
        assign out_data[1207] = lut_1207_out;
    end
    endgenerate
    
    
    
    // LUT : 1208
    wire [63:0] lut_1208_table = 64'b1100110011111101000011001100110011001100111111110000110011001100;
    wire [5:0] lut_1208_select = {
                             in_data[70],
                             in_data[345],
                             in_data[489],
                             in_data[566],
                             in_data[470],
                             in_data[306]};
    
    wire lut_1208_out = lut_1208_table[lut_1208_select];
    
    generate
    if ( USE_REG ) begin : ff_1208
        reg   lut_1208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1208_ff <= lut_1208_out;
            end
        end
        
        assign out_data[1208] = lut_1208_ff;
    end
    else begin : no_ff_1208
        assign out_data[1208] = lut_1208_out;
    end
    endgenerate
    
    
    
    // LUT : 1209
    wire [63:0] lut_1209_table = 64'b1111111111111111111111111111111111111111001010101111111100001010;
    wire [5:0] lut_1209_select = {
                             in_data[444],
                             in_data[4],
                             in_data[157],
                             in_data[409],
                             in_data[336],
                             in_data[606]};
    
    wire lut_1209_out = lut_1209_table[lut_1209_select];
    
    generate
    if ( USE_REG ) begin : ff_1209
        reg   lut_1209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1209_ff <= lut_1209_out;
            end
        end
        
        assign out_data[1209] = lut_1209_ff;
    end
    else begin : no_ff_1209
        assign out_data[1209] = lut_1209_out;
    end
    endgenerate
    
    
    
    // LUT : 1210
    wire [63:0] lut_1210_table = 64'b0101111100000000010111110000010101011111000000000101111100000101;
    wire [5:0] lut_1210_select = {
                             in_data[87],
                             in_data[777],
                             in_data[677],
                             in_data[386],
                             in_data[6],
                             in_data[106]};
    
    wire lut_1210_out = lut_1210_table[lut_1210_select];
    
    generate
    if ( USE_REG ) begin : ff_1210
        reg   lut_1210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1210_ff <= lut_1210_out;
            end
        end
        
        assign out_data[1210] = lut_1210_ff;
    end
    else begin : no_ff_1210
        assign out_data[1210] = lut_1210_out;
    end
    endgenerate
    
    
    
    // LUT : 1211
    wire [63:0] lut_1211_table = 64'b0000000000000000000000000011000000000000000100000001000000110001;
    wire [5:0] lut_1211_select = {
                             in_data[714],
                             in_data[415],
                             in_data[579],
                             in_data[598],
                             in_data[180],
                             in_data[524]};
    
    wire lut_1211_out = lut_1211_table[lut_1211_select];
    
    generate
    if ( USE_REG ) begin : ff_1211
        reg   lut_1211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1211_ff <= lut_1211_out;
            end
        end
        
        assign out_data[1211] = lut_1211_ff;
    end
    else begin : no_ff_1211
        assign out_data[1211] = lut_1211_out;
    end
    endgenerate
    
    
    
    // LUT : 1212
    wire [63:0] lut_1212_table = 64'b0101010101010101010101010101010101010101010101010101010101010101;
    wire [5:0] lut_1212_select = {
                             in_data[12],
                             in_data[173],
                             in_data[20],
                             in_data[702],
                             in_data[706],
                             in_data[403]};
    
    wire lut_1212_out = lut_1212_table[lut_1212_select];
    
    generate
    if ( USE_REG ) begin : ff_1212
        reg   lut_1212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1212_ff <= lut_1212_out;
            end
        end
        
        assign out_data[1212] = lut_1212_ff;
    end
    else begin : no_ff_1212
        assign out_data[1212] = lut_1212_out;
    end
    endgenerate
    
    
    
    // LUT : 1213
    wire [63:0] lut_1213_table = 64'b1111111100000000111111111011000011111111100000001111111111110001;
    wire [5:0] lut_1213_select = {
                             in_data[76],
                             in_data[604],
                             in_data[300],
                             in_data[188],
                             in_data[657],
                             in_data[388]};
    
    wire lut_1213_out = lut_1213_table[lut_1213_select];
    
    generate
    if ( USE_REG ) begin : ff_1213
        reg   lut_1213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1213_ff <= lut_1213_out;
            end
        end
        
        assign out_data[1213] = lut_1213_ff;
    end
    else begin : no_ff_1213
        assign out_data[1213] = lut_1213_out;
    end
    endgenerate
    
    
    
    // LUT : 1214
    wire [63:0] lut_1214_table = 64'b0101010111111111010101011111111101010101010101010101010101010101;
    wire [5:0] lut_1214_select = {
                             in_data[146],
                             in_data[731],
                             in_data[293],
                             in_data[251],
                             in_data[751],
                             in_data[408]};
    
    wire lut_1214_out = lut_1214_table[lut_1214_select];
    
    generate
    if ( USE_REG ) begin : ff_1214
        reg   lut_1214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1214_ff <= lut_1214_out;
            end
        end
        
        assign out_data[1214] = lut_1214_ff;
    end
    else begin : no_ff_1214
        assign out_data[1214] = lut_1214_out;
    end
    endgenerate
    
    
    
    // LUT : 1215
    wire [63:0] lut_1215_table = 64'b0000000011111111000100001111111100000000111111111100000011111111;
    wire [5:0] lut_1215_select = {
                             in_data[600],
                             in_data[284],
                             in_data[380],
                             in_data[561],
                             in_data[767],
                             in_data[572]};
    
    wire lut_1215_out = lut_1215_table[lut_1215_select];
    
    generate
    if ( USE_REG ) begin : ff_1215
        reg   lut_1215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1215_ff <= lut_1215_out;
            end
        end
        
        assign out_data[1215] = lut_1215_ff;
    end
    else begin : no_ff_1215
        assign out_data[1215] = lut_1215_out;
    end
    endgenerate
    
    
    
    // LUT : 1216
    wire [63:0] lut_1216_table = 64'b0111111101111111000111110000110100111111000011110001111100001100;
    wire [5:0] lut_1216_select = {
                             in_data[710],
                             in_data[243],
                             in_data[315],
                             in_data[605],
                             in_data[463],
                             in_data[552]};
    
    wire lut_1216_out = lut_1216_table[lut_1216_select];
    
    generate
    if ( USE_REG ) begin : ff_1216
        reg   lut_1216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1216_ff <= lut_1216_out;
            end
        end
        
        assign out_data[1216] = lut_1216_ff;
    end
    else begin : no_ff_1216
        assign out_data[1216] = lut_1216_out;
    end
    endgenerate
    
    
    
    // LUT : 1217
    wire [63:0] lut_1217_table = 64'b0000000100010001000001000100010000000001000100010000010001000100;
    wire [5:0] lut_1217_select = {
                             in_data[5],
                             in_data[341],
                             in_data[74],
                             in_data[724],
                             in_data[636],
                             in_data[193]};
    
    wire lut_1217_out = lut_1217_table[lut_1217_select];
    
    generate
    if ( USE_REG ) begin : ff_1217
        reg   lut_1217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1217_ff <= lut_1217_out;
            end
        end
        
        assign out_data[1217] = lut_1217_ff;
    end
    else begin : no_ff_1217
        assign out_data[1217] = lut_1217_out;
    end
    endgenerate
    
    
    
    // LUT : 1218
    wire [63:0] lut_1218_table = 64'b0101000001010100000000000101000000000000111101000010001011111111;
    wire [5:0] lut_1218_select = {
                             in_data[464],
                             in_data[407],
                             in_data[370],
                             in_data[361],
                             in_data[484],
                             in_data[317]};
    
    wire lut_1218_out = lut_1218_table[lut_1218_select];
    
    generate
    if ( USE_REG ) begin : ff_1218
        reg   lut_1218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1218_ff <= lut_1218_out;
            end
        end
        
        assign out_data[1218] = lut_1218_ff;
    end
    else begin : no_ff_1218
        assign out_data[1218] = lut_1218_out;
    end
    endgenerate
    
    
    
    // LUT : 1219
    wire [63:0] lut_1219_table = 64'b1100000011111100110000001111110011000000111111001100000011111100;
    wire [5:0] lut_1219_select = {
                             in_data[532],
                             in_data[588],
                             in_data[97],
                             in_data[658],
                             in_data[500],
                             in_data[83]};
    
    wire lut_1219_out = lut_1219_table[lut_1219_select];
    
    generate
    if ( USE_REG ) begin : ff_1219
        reg   lut_1219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1219_ff <= lut_1219_out;
            end
        end
        
        assign out_data[1219] = lut_1219_ff;
    end
    else begin : no_ff_1219
        assign out_data[1219] = lut_1219_out;
    end
    endgenerate
    
    
    
    // LUT : 1220
    wire [63:0] lut_1220_table = 64'b1100110000000000111111110000000011111111110010001111111111001110;
    wire [5:0] lut_1220_select = {
                             in_data[132],
                             in_data[770],
                             in_data[685],
                             in_data[26],
                             in_data[175],
                             in_data[757]};
    
    wire lut_1220_out = lut_1220_table[lut_1220_select];
    
    generate
    if ( USE_REG ) begin : ff_1220
        reg   lut_1220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1220_ff <= lut_1220_out;
            end
        end
        
        assign out_data[1220] = lut_1220_ff;
    end
    else begin : no_ff_1220
        assign out_data[1220] = lut_1220_out;
    end
    endgenerate
    
    
    
    // LUT : 1221
    wire [63:0] lut_1221_table = 64'b0011001111111111001100101111111100110011111111110000000000110011;
    wire [5:0] lut_1221_select = {
                             in_data[771],
                             in_data[305],
                             in_data[460],
                             in_data[504],
                             in_data[412],
                             in_data[34]};
    
    wire lut_1221_out = lut_1221_table[lut_1221_select];
    
    generate
    if ( USE_REG ) begin : ff_1221
        reg   lut_1221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1221_ff <= lut_1221_out;
            end
        end
        
        assign out_data[1221] = lut_1221_ff;
    end
    else begin : no_ff_1221
        assign out_data[1221] = lut_1221_out;
    end
    endgenerate
    
    
    
    // LUT : 1222
    wire [63:0] lut_1222_table = 64'b1110000011100000111000001111000011111000111110001110100011111100;
    wire [5:0] lut_1222_select = {
                             in_data[638],
                             in_data[138],
                             in_data[700],
                             in_data[442],
                             in_data[515],
                             in_data[462]};
    
    wire lut_1222_out = lut_1222_table[lut_1222_select];
    
    generate
    if ( USE_REG ) begin : ff_1222
        reg   lut_1222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1222_ff <= lut_1222_out;
            end
        end
        
        assign out_data[1222] = lut_1222_ff;
    end
    else begin : no_ff_1222
        assign out_data[1222] = lut_1222_out;
    end
    endgenerate
    
    
    
    // LUT : 1223
    wire [63:0] lut_1223_table = 64'b0000101010101111000011111010111100000010001011110000101000101111;
    wire [5:0] lut_1223_select = {
                             in_data[679],
                             in_data[616],
                             in_data[492],
                             in_data[181],
                             in_data[205],
                             in_data[120]};
    
    wire lut_1223_out = lut_1223_table[lut_1223_select];
    
    generate
    if ( USE_REG ) begin : ff_1223
        reg   lut_1223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1223_ff <= lut_1223_out;
            end
        end
        
        assign out_data[1223] = lut_1223_ff;
    end
    else begin : no_ff_1223
        assign out_data[1223] = lut_1223_out;
    end
    endgenerate
    
    
    
    // LUT : 1224
    wire [63:0] lut_1224_table = 64'b1010111010101010101010101010101010101010101010101010111110101010;
    wire [5:0] lut_1224_select = {
                             in_data[203],
                             in_data[601],
                             in_data[720],
                             in_data[265],
                             in_data[765],
                             in_data[482]};
    
    wire lut_1224_out = lut_1224_table[lut_1224_select];
    
    generate
    if ( USE_REG ) begin : ff_1224
        reg   lut_1224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1224_ff <= lut_1224_out;
            end
        end
        
        assign out_data[1224] = lut_1224_ff;
    end
    else begin : no_ff_1224
        assign out_data[1224] = lut_1224_out;
    end
    endgenerate
    
    
    
    // LUT : 1225
    wire [63:0] lut_1225_table = 64'b0000000011001100000000001100110000000000110011000000000011001100;
    wire [5:0] lut_1225_select = {
                             in_data[499],
                             in_data[313],
                             in_data[425],
                             in_data[255],
                             in_data[291],
                             in_data[94]};
    
    wire lut_1225_out = lut_1225_table[lut_1225_select];
    
    generate
    if ( USE_REG ) begin : ff_1225
        reg   lut_1225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1225_ff <= lut_1225_out;
            end
        end
        
        assign out_data[1225] = lut_1225_ff;
    end
    else begin : no_ff_1225
        assign out_data[1225] = lut_1225_out;
    end
    endgenerate
    
    
    
    // LUT : 1226
    wire [63:0] lut_1226_table = 64'b1100111111001100110011110000111111001111110011001110111110001111;
    wire [5:0] lut_1226_select = {
                             in_data[52],
                             in_data[508],
                             in_data[387],
                             in_data[344],
                             in_data[267],
                             in_data[773]};
    
    wire lut_1226_out = lut_1226_table[lut_1226_select];
    
    generate
    if ( USE_REG ) begin : ff_1226
        reg   lut_1226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1226_ff <= lut_1226_out;
            end
        end
        
        assign out_data[1226] = lut_1226_ff;
    end
    else begin : no_ff_1226
        assign out_data[1226] = lut_1226_out;
    end
    endgenerate
    
    
    
    // LUT : 1227
    wire [63:0] lut_1227_table = 64'b0000000010000000111111111100110011110000111100001111111111111111;
    wire [5:0] lut_1227_select = {
                             in_data[327],
                             in_data[413],
                             in_data[151],
                             in_data[369],
                             in_data[541],
                             in_data[56]};
    
    wire lut_1227_out = lut_1227_table[lut_1227_select];
    
    generate
    if ( USE_REG ) begin : ff_1227
        reg   lut_1227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1227_ff <= lut_1227_out;
            end
        end
        
        assign out_data[1227] = lut_1227_ff;
    end
    else begin : no_ff_1227
        assign out_data[1227] = lut_1227_out;
    end
    endgenerate
    
    
    
    // LUT : 1228
    wire [63:0] lut_1228_table = 64'b1111111111111111101011111110111111111111111101010000010000000000;
    wire [5:0] lut_1228_select = {
                             in_data[331],
                             in_data[343],
                             in_data[662],
                             in_data[258],
                             in_data[476],
                             in_data[509]};
    
    wire lut_1228_out = lut_1228_table[lut_1228_select];
    
    generate
    if ( USE_REG ) begin : ff_1228
        reg   lut_1228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1228_ff <= lut_1228_out;
            end
        end
        
        assign out_data[1228] = lut_1228_ff;
    end
    else begin : no_ff_1228
        assign out_data[1228] = lut_1228_out;
    end
    endgenerate
    
    
    
    // LUT : 1229
    wire [63:0] lut_1229_table = 64'b1110111111111111110011001100110011001111111011111100110011001100;
    wire [5:0] lut_1229_select = {
                             in_data[778],
                             in_data[179],
                             in_data[553],
                             in_data[268],
                             in_data[129],
                             in_data[439]};
    
    wire lut_1229_out = lut_1229_table[lut_1229_select];
    
    generate
    if ( USE_REG ) begin : ff_1229
        reg   lut_1229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1229_ff <= lut_1229_out;
            end
        end
        
        assign out_data[1229] = lut_1229_ff;
    end
    else begin : no_ff_1229
        assign out_data[1229] = lut_1229_out;
    end
    endgenerate
    
    
    
    // LUT : 1230
    wire [63:0] lut_1230_table = 64'b0101010101010101000010100000000001010101010101010000110000000000;
    wire [5:0] lut_1230_select = {
                             in_data[195],
                             in_data[514],
                             in_data[540],
                             in_data[618],
                             in_data[422],
                             in_data[426]};
    
    wire lut_1230_out = lut_1230_table[lut_1230_select];
    
    generate
    if ( USE_REG ) begin : ff_1230
        reg   lut_1230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1230_ff <= lut_1230_out;
            end
        end
        
        assign out_data[1230] = lut_1230_ff;
    end
    else begin : no_ff_1230
        assign out_data[1230] = lut_1230_out;
    end
    endgenerate
    
    
    
    // LUT : 1231
    wire [63:0] lut_1231_table = 64'b1111111100110000111111110011000111111111001100001111111100110001;
    wire [5:0] lut_1231_select = {
                             in_data[88],
                             in_data[199],
                             in_data[104],
                             in_data[332],
                             in_data[411],
                             in_data[705]};
    
    wire lut_1231_out = lut_1231_table[lut_1231_select];
    
    generate
    if ( USE_REG ) begin : ff_1231
        reg   lut_1231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1231_ff <= lut_1231_out;
            end
        end
        
        assign out_data[1231] = lut_1231_ff;
    end
    else begin : no_ff_1231
        assign out_data[1231] = lut_1231_out;
    end
    endgenerate
    
    
    
    // LUT : 1232
    wire [63:0] lut_1232_table = 64'b0000000000000010000000100000111100000000000000000000000000001000;
    wire [5:0] lut_1232_select = {
                             in_data[545],
                             in_data[633],
                             in_data[594],
                             in_data[635],
                             in_data[136],
                             in_data[431]};
    
    wire lut_1232_out = lut_1232_table[lut_1232_select];
    
    generate
    if ( USE_REG ) begin : ff_1232
        reg   lut_1232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1232_ff <= lut_1232_out;
            end
        end
        
        assign out_data[1232] = lut_1232_ff;
    end
    else begin : no_ff_1232
        assign out_data[1232] = lut_1232_out;
    end
    endgenerate
    
    
    
    // LUT : 1233
    wire [63:0] lut_1233_table = 64'b0011011100000000111111110000000000000000000000000000000100000000;
    wire [5:0] lut_1233_select = {
                             in_data[519],
                             in_data[626],
                             in_data[465],
                             in_data[137],
                             in_data[190],
                             in_data[22]};
    
    wire lut_1233_out = lut_1233_table[lut_1233_select];
    
    generate
    if ( USE_REG ) begin : ff_1233
        reg   lut_1233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1233_ff <= lut_1233_out;
            end
        end
        
        assign out_data[1233] = lut_1233_ff;
    end
    else begin : no_ff_1233
        assign out_data[1233] = lut_1233_out;
    end
    endgenerate
    
    
    
    // LUT : 1234
    wire [63:0] lut_1234_table = 64'b1111010111111111010101011111111100000000000000000000000000000000;
    wire [5:0] lut_1234_select = {
                             in_data[347],
                             in_data[473],
                             in_data[290],
                             in_data[617],
                             in_data[338],
                             in_data[440]};
    
    wire lut_1234_out = lut_1234_table[lut_1234_select];
    
    generate
    if ( USE_REG ) begin : ff_1234
        reg   lut_1234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1234_ff <= lut_1234_out;
            end
        end
        
        assign out_data[1234] = lut_1234_ff;
    end
    else begin : no_ff_1234
        assign out_data[1234] = lut_1234_out;
    end
    endgenerate
    
    
    
    // LUT : 1235
    wire [63:0] lut_1235_table = 64'b0000000100000001000000010000000100000000000000010000000100000001;
    wire [5:0] lut_1235_select = {
                             in_data[764],
                             in_data[152],
                             in_data[446],
                             in_data[659],
                             in_data[608],
                             in_data[330]};
    
    wire lut_1235_out = lut_1235_table[lut_1235_select];
    
    generate
    if ( USE_REG ) begin : ff_1235
        reg   lut_1235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1235_ff <= lut_1235_out;
            end
        end
        
        assign out_data[1235] = lut_1235_ff;
    end
    else begin : no_ff_1235
        assign out_data[1235] = lut_1235_out;
    end
    endgenerate
    
    
    
    // LUT : 1236
    wire [63:0] lut_1236_table = 64'b1100110111001101110011001100110011001100110011011100110011001100;
    wire [5:0] lut_1236_select = {
                             in_data[61],
                             in_data[754],
                             in_data[60],
                             in_data[350],
                             in_data[234],
                             in_data[122]};
    
    wire lut_1236_out = lut_1236_table[lut_1236_select];
    
    generate
    if ( USE_REG ) begin : ff_1236
        reg   lut_1236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1236_ff <= lut_1236_out;
            end
        end
        
        assign out_data[1236] = lut_1236_ff;
    end
    else begin : no_ff_1236
        assign out_data[1236] = lut_1236_out;
    end
    endgenerate
    
    
    
    // LUT : 1237
    wire [63:0] lut_1237_table = 64'b1111000011111010111111101111111101000000111110101110100011111110;
    wire [5:0] lut_1237_select = {
                             in_data[454],
                             in_data[379],
                             in_data[708],
                             in_data[637],
                             in_data[595],
                             in_data[399]};
    
    wire lut_1237_out = lut_1237_table[lut_1237_select];
    
    generate
    if ( USE_REG ) begin : ff_1237
        reg   lut_1237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1237_ff <= lut_1237_out;
            end
        end
        
        assign out_data[1237] = lut_1237_ff;
    end
    else begin : no_ff_1237
        assign out_data[1237] = lut_1237_out;
    end
    endgenerate
    
    
    
    // LUT : 1238
    wire [63:0] lut_1238_table = 64'b0000000000000000010100110101011100000000000000000101001100010011;
    wire [5:0] lut_1238_select = {
                             in_data[7],
                             in_data[185],
                             in_data[762],
                             in_data[577],
                             in_data[150],
                             in_data[619]};
    
    wire lut_1238_out = lut_1238_table[lut_1238_select];
    
    generate
    if ( USE_REG ) begin : ff_1238
        reg   lut_1238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1238_ff <= lut_1238_out;
            end
        end
        
        assign out_data[1238] = lut_1238_ff;
    end
    else begin : no_ff_1238
        assign out_data[1238] = lut_1238_out;
    end
    endgenerate
    
    
    
    // LUT : 1239
    wire [63:0] lut_1239_table = 64'b1101010111010101110101011111010101000000010000000101000001010000;
    wire [5:0] lut_1239_select = {
                             in_data[493],
                             in_data[335],
                             in_data[421],
                             in_data[42],
                             in_data[779],
                             in_data[390]};
    
    wire lut_1239_out = lut_1239_table[lut_1239_select];
    
    generate
    if ( USE_REG ) begin : ff_1239
        reg   lut_1239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1239_ff <= lut_1239_out;
            end
        end
        
        assign out_data[1239] = lut_1239_ff;
    end
    else begin : no_ff_1239
        assign out_data[1239] = lut_1239_out;
    end
    endgenerate
    
    
    
    // LUT : 1240
    wire [63:0] lut_1240_table = 64'b1110111111101111010011110100111100001000000010000000000000000000;
    wire [5:0] lut_1240_select = {
                             in_data[466],
                             in_data[264],
                             in_data[92],
                             in_data[689],
                             in_data[653],
                             in_data[438]};
    
    wire lut_1240_out = lut_1240_table[lut_1240_select];
    
    generate
    if ( USE_REG ) begin : ff_1240
        reg   lut_1240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1240_ff <= lut_1240_out;
            end
        end
        
        assign out_data[1240] = lut_1240_ff;
    end
    else begin : no_ff_1240
        assign out_data[1240] = lut_1240_out;
    end
    endgenerate
    
    
    
    // LUT : 1241
    wire [63:0] lut_1241_table = 64'b0000111111111111000000001111111100001111111111110000111101001111;
    wire [5:0] lut_1241_select = {
                             in_data[204],
                             in_data[339],
                             in_data[215],
                             in_data[208],
                             in_data[15],
                             in_data[506]};
    
    wire lut_1241_out = lut_1241_table[lut_1241_select];
    
    generate
    if ( USE_REG ) begin : ff_1241
        reg   lut_1241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1241_ff <= lut_1241_out;
            end
        end
        
        assign out_data[1241] = lut_1241_ff;
    end
    else begin : no_ff_1241
        assign out_data[1241] = lut_1241_out;
    end
    endgenerate
    
    
    
    // LUT : 1242
    wire [63:0] lut_1242_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_1242_select = {
                             in_data[397],
                             in_data[551],
                             in_data[656],
                             in_data[477],
                             in_data[450],
                             in_data[367]};
    
    wire lut_1242_out = lut_1242_table[lut_1242_select];
    
    generate
    if ( USE_REG ) begin : ff_1242
        reg   lut_1242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1242_ff <= lut_1242_out;
            end
        end
        
        assign out_data[1242] = lut_1242_ff;
    end
    else begin : no_ff_1242
        assign out_data[1242] = lut_1242_out;
    end
    endgenerate
    
    
    
    // LUT : 1243
    wire [63:0] lut_1243_table = 64'b1111000011110000111111001111000011111110111100001111111111110000;
    wire [5:0] lut_1243_select = {
                             in_data[452],
                             in_data[494],
                             in_data[322],
                             in_data[155],
                             in_data[417],
                             in_data[8]};
    
    wire lut_1243_out = lut_1243_table[lut_1243_select];
    
    generate
    if ( USE_REG ) begin : ff_1243
        reg   lut_1243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1243_ff <= lut_1243_out;
            end
        end
        
        assign out_data[1243] = lut_1243_ff;
    end
    else begin : no_ff_1243
        assign out_data[1243] = lut_1243_out;
    end
    endgenerate
    
    
    
    // LUT : 1244
    wire [63:0] lut_1244_table = 64'b1111111111111111111100001111110011111011111111111111000011111000;
    wire [5:0] lut_1244_select = {
                             in_data[364],
                             in_data[526],
                             in_data[321],
                             in_data[661],
                             in_data[99],
                             in_data[21]};
    
    wire lut_1244_out = lut_1244_table[lut_1244_select];
    
    generate
    if ( USE_REG ) begin : ff_1244
        reg   lut_1244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1244_ff <= lut_1244_out;
            end
        end
        
        assign out_data[1244] = lut_1244_ff;
    end
    else begin : no_ff_1244
        assign out_data[1244] = lut_1244_out;
    end
    endgenerate
    
    
    
    // LUT : 1245
    wire [63:0] lut_1245_table = 64'b0000000000000001000000000001010100000000000000010000000000010101;
    wire [5:0] lut_1245_select = {
                             in_data[730],
                             in_data[118],
                             in_data[124],
                             in_data[627],
                             in_data[348],
                             in_data[218]};
    
    wire lut_1245_out = lut_1245_table[lut_1245_select];
    
    generate
    if ( USE_REG ) begin : ff_1245
        reg   lut_1245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1245_ff <= lut_1245_out;
            end
        end
        
        assign out_data[1245] = lut_1245_ff;
    end
    else begin : no_ff_1245
        assign out_data[1245] = lut_1245_out;
    end
    endgenerate
    
    
    
    // LUT : 1246
    wire [63:0] lut_1246_table = 64'b0000100000000000111111110000110011111111000000111111111100110111;
    wire [5:0] lut_1246_select = {
                             in_data[435],
                             in_data[517],
                             in_data[383],
                             in_data[66],
                             in_data[544],
                             in_data[759]};
    
    wire lut_1246_out = lut_1246_table[lut_1246_select];
    
    generate
    if ( USE_REG ) begin : ff_1246
        reg   lut_1246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1246_ff <= lut_1246_out;
            end
        end
        
        assign out_data[1246] = lut_1246_ff;
    end
    else begin : no_ff_1246
        assign out_data[1246] = lut_1246_out;
    end
    endgenerate
    
    
    
    // LUT : 1247
    wire [63:0] lut_1247_table = 64'b1111111100000000111111111000110011111111110011001111111111001100;
    wire [5:0] lut_1247_select = {
                             in_data[183],
                             in_data[480],
                             in_data[192],
                             in_data[563],
                             in_data[602],
                             in_data[394]};
    
    wire lut_1247_out = lut_1247_table[lut_1247_select];
    
    generate
    if ( USE_REG ) begin : ff_1247
        reg   lut_1247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1247_ff <= lut_1247_out;
            end
        end
        
        assign out_data[1247] = lut_1247_ff;
    end
    else begin : no_ff_1247
        assign out_data[1247] = lut_1247_out;
    end
    endgenerate
    
    
    
    // LUT : 1248
    wire [63:0] lut_1248_table = 64'b0000111100001111000011110000111100001111000011110000111100001111;
    wire [5:0] lut_1248_select = {
                             in_data[311],
                             in_data[647],
                             in_data[782],
                             in_data[488],
                             in_data[48],
                             in_data[170]};
    
    wire lut_1248_out = lut_1248_table[lut_1248_select];
    
    generate
    if ( USE_REG ) begin : ff_1248
        reg   lut_1248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1248_ff <= lut_1248_out;
            end
        end
        
        assign out_data[1248] = lut_1248_ff;
    end
    else begin : no_ff_1248
        assign out_data[1248] = lut_1248_out;
    end
    endgenerate
    
    
    
    // LUT : 1249
    wire [63:0] lut_1249_table = 64'b0111000000110000011100000011000011110000011100001111010111110000;
    wire [5:0] lut_1249_select = {
                             in_data[351],
                             in_data[277],
                             in_data[172],
                             in_data[398],
                             in_data[622],
                             in_data[72]};
    
    wire lut_1249_out = lut_1249_table[lut_1249_select];
    
    generate
    if ( USE_REG ) begin : ff_1249
        reg   lut_1249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1249_ff <= lut_1249_out;
            end
        end
        
        assign out_data[1249] = lut_1249_ff;
    end
    else begin : no_ff_1249
        assign out_data[1249] = lut_1249_out;
    end
    endgenerate
    
    
    
    // LUT : 1250
    wire [63:0] lut_1250_table = 64'b0111011101110111010101010101010101110111010101010101010101010101;
    wire [5:0] lut_1250_select = {
                             in_data[557],
                             in_data[581],
                             in_data[590],
                             in_data[531],
                             in_data[275],
                             in_data[542]};
    
    wire lut_1250_out = lut_1250_table[lut_1250_select];
    
    generate
    if ( USE_REG ) begin : ff_1250
        reg   lut_1250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1250_ff <= lut_1250_out;
            end
        end
        
        assign out_data[1250] = lut_1250_ff;
    end
    else begin : no_ff_1250
        assign out_data[1250] = lut_1250_out;
    end
    endgenerate
    
    
    
    // LUT : 1251
    wire [63:0] lut_1251_table = 64'b1110111011111111111111111111111111101110111011101010101011101110;
    wire [5:0] lut_1251_select = {
                             in_data[678],
                             in_data[377],
                             in_data[147],
                             in_data[89],
                             in_data[660],
                             in_data[274]};
    
    wire lut_1251_out = lut_1251_table[lut_1251_select];
    
    generate
    if ( USE_REG ) begin : ff_1251
        reg   lut_1251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1251_ff <= lut_1251_out;
            end
        end
        
        assign out_data[1251] = lut_1251_ff;
    end
    else begin : no_ff_1251
        assign out_data[1251] = lut_1251_out;
    end
    endgenerate
    
    
    
    // LUT : 1252
    wire [63:0] lut_1252_table = 64'b0111010101110100011101000111010001110100011101000111010001110100;
    wire [5:0] lut_1252_select = {
                             in_data[119],
                             in_data[135],
                             in_data[25],
                             in_data[156],
                             in_data[432],
                             in_data[304]};
    
    wire lut_1252_out = lut_1252_table[lut_1252_select];
    
    generate
    if ( USE_REG ) begin : ff_1252
        reg   lut_1252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1252_ff <= lut_1252_out;
            end
        end
        
        assign out_data[1252] = lut_1252_ff;
    end
    else begin : no_ff_1252
        assign out_data[1252] = lut_1252_out;
    end
    endgenerate
    
    
    
    // LUT : 1253
    wire [63:0] lut_1253_table = 64'b1111111111111111111111111111111101000101000001000000010000000000;
    wire [5:0] lut_1253_select = {
                             in_data[603],
                             in_data[178],
                             in_data[501],
                             in_data[613],
                             in_data[78],
                             in_data[640]};
    
    wire lut_1253_out = lut_1253_table[lut_1253_select];
    
    generate
    if ( USE_REG ) begin : ff_1253
        reg   lut_1253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1253_ff <= lut_1253_out;
            end
        end
        
        assign out_data[1253] = lut_1253_ff;
    end
    else begin : no_ff_1253
        assign out_data[1253] = lut_1253_out;
    end
    endgenerate
    
    
    
    // LUT : 1254
    wire [63:0] lut_1254_table = 64'b0000000000000100000000000000000000001111000011110000111100000000;
    wire [5:0] lut_1254_select = {
                             in_data[461],
                             in_data[575],
                             in_data[510],
                             in_data[688],
                             in_data[363],
                             in_data[744]};
    
    wire lut_1254_out = lut_1254_table[lut_1254_select];
    
    generate
    if ( USE_REG ) begin : ff_1254
        reg   lut_1254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1254_ff <= lut_1254_out;
            end
        end
        
        assign out_data[1254] = lut_1254_ff;
    end
    else begin : no_ff_1254
        assign out_data[1254] = lut_1254_out;
    end
    endgenerate
    
    
    
    // LUT : 1255
    wire [63:0] lut_1255_table = 64'b0000000000000000010101010000000000000000000000000101010100000000;
    wire [5:0] lut_1255_select = {
                             in_data[169],
                             in_data[230],
                             in_data[574],
                             in_data[210],
                             in_data[211],
                             in_data[681]};
    
    wire lut_1255_out = lut_1255_table[lut_1255_select];
    
    generate
    if ( USE_REG ) begin : ff_1255
        reg   lut_1255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1255_ff <= lut_1255_out;
            end
        end
        
        assign out_data[1255] = lut_1255_ff;
    end
    else begin : no_ff_1255
        assign out_data[1255] = lut_1255_out;
    end
    endgenerate
    
    
    
    // LUT : 1256
    wire [63:0] lut_1256_table = 64'b0000000000000000001100110011001100000000000000000011001100110011;
    wire [5:0] lut_1256_select = {
                             in_data[141],
                             in_data[79],
                             in_data[45],
                             in_data[86],
                             in_data[239],
                             in_data[448]};
    
    wire lut_1256_out = lut_1256_table[lut_1256_select];
    
    generate
    if ( USE_REG ) begin : ff_1256
        reg   lut_1256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1256_ff <= lut_1256_out;
            end
        end
        
        assign out_data[1256] = lut_1256_ff;
    end
    else begin : no_ff_1256
        assign out_data[1256] = lut_1256_out;
    end
    endgenerate
    
    
    
    // LUT : 1257
    wire [63:0] lut_1257_table = 64'b0000000001000100010001001100110000000000110011000100010011011101;
    wire [5:0] lut_1257_select = {
                             in_data[247],
                             in_data[580],
                             in_data[666],
                             in_data[587],
                             in_data[164],
                             in_data[745]};
    
    wire lut_1257_out = lut_1257_table[lut_1257_select];
    
    generate
    if ( USE_REG ) begin : ff_1257
        reg   lut_1257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1257_ff <= lut_1257_out;
            end
        end
        
        assign out_data[1257] = lut_1257_ff;
    end
    else begin : no_ff_1257
        assign out_data[1257] = lut_1257_out;
    end
    endgenerate
    
    
    
    // LUT : 1258
    wire [63:0] lut_1258_table = 64'b1101010011010100110101001101010011111111111111111111110011111100;
    wire [5:0] lut_1258_select = {
                             in_data[548],
                             in_data[690],
                             in_data[783],
                             in_data[214],
                             in_data[340],
                             in_data[591]};
    
    wire lut_1258_out = lut_1258_table[lut_1258_select];
    
    generate
    if ( USE_REG ) begin : ff_1258
        reg   lut_1258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1258_ff <= lut_1258_out;
            end
        end
        
        assign out_data[1258] = lut_1258_ff;
    end
    else begin : no_ff_1258
        assign out_data[1258] = lut_1258_out;
    end
    endgenerate
    
    
    
    // LUT : 1259
    wire [63:0] lut_1259_table = 64'b1100010011111111111111111100110000000000010011001111111111111100;
    wire [5:0] lut_1259_select = {
                             in_data[288],
                             in_data[154],
                             in_data[596],
                             in_data[537],
                             in_data[362],
                             in_data[768]};
    
    wire lut_1259_out = lut_1259_table[lut_1259_select];
    
    generate
    if ( USE_REG ) begin : ff_1259
        reg   lut_1259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1259_ff <= lut_1259_out;
            end
        end
        
        assign out_data[1259] = lut_1259_ff;
    end
    else begin : no_ff_1259
        assign out_data[1259] = lut_1259_out;
    end
    endgenerate
    
    
    
    // LUT : 1260
    wire [63:0] lut_1260_table = 64'b1111111110101010101010101010101011111111111111111111111110101010;
    wire [5:0] lut_1260_select = {
                             in_data[676],
                             in_data[37],
                             in_data[682],
                             in_data[28],
                             in_data[672],
                             in_data[535]};
    
    wire lut_1260_out = lut_1260_table[lut_1260_select];
    
    generate
    if ( USE_REG ) begin : ff_1260
        reg   lut_1260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1260_ff <= lut_1260_out;
            end
        end
        
        assign out_data[1260] = lut_1260_ff;
    end
    else begin : no_ff_1260
        assign out_data[1260] = lut_1260_out;
    end
    endgenerate
    
    
    
    // LUT : 1261
    wire [63:0] lut_1261_table = 64'b1111000011111100110100001111000011111100111111001100000011001000;
    wire [5:0] lut_1261_select = {
                             in_data[270],
                             in_data[316],
                             in_data[663],
                             in_data[428],
                             in_data[400],
                             in_data[140]};
    
    wire lut_1261_out = lut_1261_table[lut_1261_select];
    
    generate
    if ( USE_REG ) begin : ff_1261
        reg   lut_1261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1261_ff <= lut_1261_out;
            end
        end
        
        assign out_data[1261] = lut_1261_ff;
    end
    else begin : no_ff_1261
        assign out_data[1261] = lut_1261_out;
    end
    endgenerate
    
    
    
    // LUT : 1262
    wire [63:0] lut_1262_table = 64'b0000000010111011000000001011111100000000100010000000000010111011;
    wire [5:0] lut_1262_select = {
                             in_data[334],
                             in_data[187],
                             in_data[652],
                             in_data[82],
                             in_data[148],
                             in_data[522]};
    
    wire lut_1262_out = lut_1262_table[lut_1262_select];
    
    generate
    if ( USE_REG ) begin : ff_1262
        reg   lut_1262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1262_ff <= lut_1262_out;
            end
        end
        
        assign out_data[1262] = lut_1262_ff;
    end
    else begin : no_ff_1262
        assign out_data[1262] = lut_1262_out;
    end
    endgenerate
    
    
    
    // LUT : 1263
    wire [63:0] lut_1263_table = 64'b1111111111111111111111111111111111111111111111110000000000001010;
    wire [5:0] lut_1263_select = {
                             in_data[534],
                             in_data[649],
                             in_data[279],
                             in_data[420],
                             in_data[224],
                             in_data[696]};
    
    wire lut_1263_out = lut_1263_table[lut_1263_select];
    
    generate
    if ( USE_REG ) begin : ff_1263
        reg   lut_1263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1263_ff <= lut_1263_out;
            end
        end
        
        assign out_data[1263] = lut_1263_ff;
    end
    else begin : no_ff_1263
        assign out_data[1263] = lut_1263_out;
    end
    endgenerate
    
    
    
    // LUT : 1264
    wire [63:0] lut_1264_table = 64'b0000000000000000000000000000000000000000000000000000000011111111;
    wire [5:0] lut_1264_select = {
                             in_data[402],
                             in_data[747],
                             in_data[732],
                             in_data[13],
                             in_data[57],
                             in_data[36]};
    
    wire lut_1264_out = lut_1264_table[lut_1264_select];
    
    generate
    if ( USE_REG ) begin : ff_1264
        reg   lut_1264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1264_ff <= lut_1264_out;
            end
        end
        
        assign out_data[1264] = lut_1264_ff;
    end
    else begin : no_ff_1264
        assign out_data[1264] = lut_1264_out;
    end
    endgenerate
    
    
    
    // LUT : 1265
    wire [63:0] lut_1265_table = 64'b0000000000000000111111111111111100000000000000001111111111111111;
    wire [5:0] lut_1265_select = {
                             in_data[774],
                             in_data[217],
                             in_data[404],
                             in_data[168],
                             in_data[91],
                             in_data[673]};
    
    wire lut_1265_out = lut_1265_table[lut_1265_select];
    
    generate
    if ( USE_REG ) begin : ff_1265
        reg   lut_1265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1265_ff <= lut_1265_out;
            end
        end
        
        assign out_data[1265] = lut_1265_ff;
    end
    else begin : no_ff_1265
        assign out_data[1265] = lut_1265_out;
    end
    endgenerate
    
    
    
    // LUT : 1266
    wire [63:0] lut_1266_table = 64'b1111101111110001111100111111000011111111111100011111001111110000;
    wire [5:0] lut_1266_select = {
                             in_data[281],
                             in_data[144],
                             in_data[451],
                             in_data[299],
                             in_data[209],
                             in_data[54]};
    
    wire lut_1266_out = lut_1266_table[lut_1266_select];
    
    generate
    if ( USE_REG ) begin : ff_1266
        reg   lut_1266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1266_ff <= lut_1266_out;
            end
        end
        
        assign out_data[1266] = lut_1266_ff;
    end
    else begin : no_ff_1266
        assign out_data[1266] = lut_1266_out;
    end
    endgenerate
    
    
    
    // LUT : 1267
    wire [63:0] lut_1267_table = 64'b1010001010100000101010111010101010100010101000001011101110101010;
    wire [5:0] lut_1267_select = {
                             in_data[41],
                             in_data[564],
                             in_data[641],
                             in_data[244],
                             in_data[254],
                             in_data[358]};
    
    wire lut_1267_out = lut_1267_table[lut_1267_select];
    
    generate
    if ( USE_REG ) begin : ff_1267
        reg   lut_1267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1267_ff <= lut_1267_out;
            end
        end
        
        assign out_data[1267] = lut_1267_ff;
    end
    else begin : no_ff_1267
        assign out_data[1267] = lut_1267_out;
    end
    endgenerate
    
    
    
    // LUT : 1268
    wire [63:0] lut_1268_table = 64'b1110000011111010111000001111101010100000111110001010000011111010;
    wire [5:0] lut_1268_select = {
                             in_data[47],
                             in_data[225],
                             in_data[312],
                             in_data[406],
                             in_data[728],
                             in_data[623]};
    
    wire lut_1268_out = lut_1268_table[lut_1268_select];
    
    generate
    if ( USE_REG ) begin : ff_1268
        reg   lut_1268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1268_ff <= lut_1268_out;
            end
        end
        
        assign out_data[1268] = lut_1268_ff;
    end
    else begin : no_ff_1268
        assign out_data[1268] = lut_1268_out;
    end
    endgenerate
    
    
    
    // LUT : 1269
    wire [63:0] lut_1269_table = 64'b0101110111111101000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1269_select = {
                             in_data[233],
                             in_data[474],
                             in_data[19],
                             in_data[1],
                             in_data[252],
                             in_data[755]};
    
    wire lut_1269_out = lut_1269_table[lut_1269_select];
    
    generate
    if ( USE_REG ) begin : ff_1269
        reg   lut_1269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1269_ff <= lut_1269_out;
            end
        end
        
        assign out_data[1269] = lut_1269_ff;
    end
    else begin : no_ff_1269
        assign out_data[1269] = lut_1269_out;
    end
    endgenerate
    
    
    
    // LUT : 1270
    wire [63:0] lut_1270_table = 64'b1111111111111111111111111111000011111111111111111111111111110000;
    wire [5:0] lut_1270_select = {
                             in_data[750],
                             in_data[276],
                             in_data[376],
                             in_data[158],
                             in_data[53],
                             in_data[10]};
    
    wire lut_1270_out = lut_1270_table[lut_1270_select];
    
    generate
    if ( USE_REG ) begin : ff_1270
        reg   lut_1270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1270_ff <= lut_1270_out;
            end
        end
        
        assign out_data[1270] = lut_1270_ff;
    end
    else begin : no_ff_1270
        assign out_data[1270] = lut_1270_out;
    end
    endgenerate
    
    
    
    // LUT : 1271
    wire [63:0] lut_1271_table = 64'b0000111100000000111111110000100011101111000000001111111100001111;
    wire [5:0] lut_1271_select = {
                             in_data[625],
                             in_data[326],
                             in_data[121],
                             in_data[220],
                             in_data[112],
                             in_data[282]};
    
    wire lut_1271_out = lut_1271_table[lut_1271_select];
    
    generate
    if ( USE_REG ) begin : ff_1271
        reg   lut_1271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1271_ff <= lut_1271_out;
            end
        end
        
        assign out_data[1271] = lut_1271_ff;
    end
    else begin : no_ff_1271
        assign out_data[1271] = lut_1271_out;
    end
    endgenerate
    
    
    
    // LUT : 1272
    wire [63:0] lut_1272_table = 64'b0001000100010001110111011111111100000000000000001101110111011101;
    wire [5:0] lut_1272_select = {
                             in_data[371],
                             in_data[495],
                             in_data[165],
                             in_data[775],
                             in_data[607],
                             in_data[686]};
    
    wire lut_1272_out = lut_1272_table[lut_1272_select];
    
    generate
    if ( USE_REG ) begin : ff_1272
        reg   lut_1272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1272_ff <= lut_1272_out;
            end
        end
        
        assign out_data[1272] = lut_1272_ff;
    end
    else begin : no_ff_1272
        assign out_data[1272] = lut_1272_out;
    end
    endgenerate
    
    
    
    // LUT : 1273
    wire [63:0] lut_1273_table = 64'b1100110010000000111111111100110011001100110011001111111111011100;
    wire [5:0] lut_1273_select = {
                             in_data[44],
                             in_data[453],
                             in_data[443],
                             in_data[64],
                             in_data[126],
                             in_data[781]};
    
    wire lut_1273_out = lut_1273_table[lut_1273_select];
    
    generate
    if ( USE_REG ) begin : ff_1273
        reg   lut_1273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1273_ff <= lut_1273_out;
            end
        end
        
        assign out_data[1273] = lut_1273_ff;
    end
    else begin : no_ff_1273
        assign out_data[1273] = lut_1273_out;
    end
    endgenerate
    
    
    
    // LUT : 1274
    wire [63:0] lut_1274_table = 64'b1111101110101010111110111110110011111011101010101111101111101100;
    wire [5:0] lut_1274_select = {
                             in_data[143],
                             in_data[485],
                             in_data[543],
                             in_data[80],
                             in_data[271],
                             in_data[716]};
    
    wire lut_1274_out = lut_1274_table[lut_1274_select];
    
    generate
    if ( USE_REG ) begin : ff_1274
        reg   lut_1274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1274_ff <= lut_1274_out;
            end
        end
        
        assign out_data[1274] = lut_1274_ff;
    end
    else begin : no_ff_1274
        assign out_data[1274] = lut_1274_out;
    end
    endgenerate
    
    
    
    // LUT : 1275
    wire [63:0] lut_1275_table = 64'b1111111111111111111111111011111111111111111111111111111100000000;
    wire [5:0] lut_1275_select = {
                             in_data[693],
                             in_data[184],
                             in_data[513],
                             in_data[310],
                             in_data[475],
                             in_data[503]};
    
    wire lut_1275_out = lut_1275_table[lut_1275_select];
    
    generate
    if ( USE_REG ) begin : ff_1275
        reg   lut_1275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1275_ff <= lut_1275_out;
            end
        end
        
        assign out_data[1275] = lut_1275_ff;
    end
    else begin : no_ff_1275
        assign out_data[1275] = lut_1275_out;
    end
    endgenerate
    
    
    
    // LUT : 1276
    wire [63:0] lut_1276_table = 64'b1100110011001100000000000000000011111110110011000011001100110011;
    wire [5:0] lut_1276_select = {
                             in_data[65],
                             in_data[573],
                             in_data[392],
                             in_data[725],
                             in_data[683],
                             in_data[9]};
    
    wire lut_1276_out = lut_1276_table[lut_1276_select];
    
    generate
    if ( USE_REG ) begin : ff_1276
        reg   lut_1276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1276_ff <= lut_1276_out;
            end
        end
        
        assign out_data[1276] = lut_1276_ff;
    end
    else begin : no_ff_1276
        assign out_data[1276] = lut_1276_out;
    end
    endgenerate
    
    
    
    // LUT : 1277
    wire [63:0] lut_1277_table = 64'b1011111111111111101010101010101011111111111111111111111111111111;
    wire [5:0] lut_1277_select = {
                             in_data[206],
                             in_data[162],
                             in_data[31],
                             in_data[63],
                             in_data[447],
                             in_data[159]};
    
    wire lut_1277_out = lut_1277_table[lut_1277_select];
    
    generate
    if ( USE_REG ) begin : ff_1277
        reg   lut_1277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1277_ff <= lut_1277_out;
            end
        end
        
        assign out_data[1277] = lut_1277_ff;
    end
    else begin : no_ff_1277
        assign out_data[1277] = lut_1277_out;
    end
    endgenerate
    
    
    
    // LUT : 1278
    wire [63:0] lut_1278_table = 64'b1110111110101111111011111010111111111111101011111110111100101111;
    wire [5:0] lut_1278_select = {
                             in_data[760],
                             in_data[73],
                             in_data[718],
                             in_data[523],
                             in_data[739],
                             in_data[630]};
    
    wire lut_1278_out = lut_1278_table[lut_1278_select];
    
    generate
    if ( USE_REG ) begin : ff_1278
        reg   lut_1278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1278_ff <= lut_1278_out;
            end
        end
        
        assign out_data[1278] = lut_1278_ff;
    end
    else begin : no_ff_1278
        assign out_data[1278] = lut_1278_out;
    end
    endgenerate
    
    
    
    // LUT : 1279
    wire [63:0] lut_1279_table = 64'b1111111111111111111111111111111111111101111111001111110011111100;
    wire [5:0] lut_1279_select = {
                             in_data[95],
                             in_data[772],
                             in_data[43],
                             in_data[502],
                             in_data[550],
                             in_data[116]};
    
    wire lut_1279_out = lut_1279_table[lut_1279_select];
    
    generate
    if ( USE_REG ) begin : ff_1279
        reg   lut_1279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1279_ff <= lut_1279_out;
            end
        end
        
        assign out_data[1279] = lut_1279_ff;
    end
    else begin : no_ff_1279
        assign out_data[1279] = lut_1279_out;
    end
    endgenerate
    
    
    
    // LUT : 1280
    wire [63:0] lut_1280_table = 64'b0100111100001111000000000000101111111010000011111000101000001111;
    wire [5:0] lut_1280_select = {
                             in_data[130],
                             in_data[71],
                             in_data[437],
                             in_data[352],
                             in_data[669],
                             in_data[235]};
    
    wire lut_1280_out = lut_1280_table[lut_1280_select];
    
    generate
    if ( USE_REG ) begin : ff_1280
        reg   lut_1280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1280_ff <= lut_1280_out;
            end
        end
        
        assign out_data[1280] = lut_1280_ff;
    end
    else begin : no_ff_1280
        assign out_data[1280] = lut_1280_out;
    end
    endgenerate
    
    
    
    // LUT : 1281
    wire [63:0] lut_1281_table = 64'b1111111111111111111111111111111111111111000101011111111100000000;
    wire [5:0] lut_1281_select = {
                             in_data[257],
                             in_data[472],
                             in_data[216],
                             in_data[226],
                             in_data[337],
                             in_data[478]};
    
    wire lut_1281_out = lut_1281_table[lut_1281_select];
    
    generate
    if ( USE_REG ) begin : ff_1281
        reg   lut_1281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1281_ff <= lut_1281_out;
            end
        end
        
        assign out_data[1281] = lut_1281_ff;
    end
    else begin : no_ff_1281
        assign out_data[1281] = lut_1281_out;
    end
    endgenerate
    
    
    
    // LUT : 1282
    wire [63:0] lut_1282_table = 64'b1111111111111111101011111010101011111111111111111010111110101011;
    wire [5:0] lut_1282_select = {
                             in_data[280],
                             in_data[131],
                             in_data[256],
                             in_data[546],
                             in_data[110],
                             in_data[684]};
    
    wire lut_1282_out = lut_1282_table[lut_1282_select];
    
    generate
    if ( USE_REG ) begin : ff_1282
        reg   lut_1282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1282_ff <= lut_1282_out;
            end
        end
        
        assign out_data[1282] = lut_1282_ff;
    end
    else begin : no_ff_1282
        assign out_data[1282] = lut_1282_out;
    end
    endgenerate
    
    
    
    // LUT : 1283
    wire [63:0] lut_1283_table = 64'b1111111111110000111100001111000011111111111100001111000011110000;
    wire [5:0] lut_1283_select = {
                             in_data[16],
                             in_data[721],
                             in_data[490],
                             in_data[318],
                             in_data[23],
                             in_data[14]};
    
    wire lut_1283_out = lut_1283_table[lut_1283_select];
    
    generate
    if ( USE_REG ) begin : ff_1283
        reg   lut_1283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1283_ff <= lut_1283_out;
            end
        end
        
        assign out_data[1283] = lut_1283_ff;
    end
    else begin : no_ff_1283
        assign out_data[1283] = lut_1283_out;
    end
    endgenerate
    
    
    
    // LUT : 1284
    wire [63:0] lut_1284_table = 64'b1111111111111111000011000000000011111111111111110000110000000100;
    wire [5:0] lut_1284_select = {
                             in_data[756],
                             in_data[459],
                             in_data[85],
                             in_data[96],
                             in_data[103],
                             in_data[670]};
    
    wire lut_1284_out = lut_1284_table[lut_1284_select];
    
    generate
    if ( USE_REG ) begin : ff_1284
        reg   lut_1284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1284_ff <= lut_1284_out;
            end
        end
        
        assign out_data[1284] = lut_1284_ff;
    end
    else begin : no_ff_1284
        assign out_data[1284] = lut_1284_out;
    end
    endgenerate
    
    
    
    // LUT : 1285
    wire [63:0] lut_1285_table = 64'b1111111100000101010111110000010111111111000001000101111100000000;
    wire [5:0] lut_1285_select = {
                             in_data[445],
                             in_data[483],
                             in_data[349],
                             in_data[289],
                             in_data[559],
                             in_data[145]};
    
    wire lut_1285_out = lut_1285_table[lut_1285_select];
    
    generate
    if ( USE_REG ) begin : ff_1285
        reg   lut_1285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1285_ff <= lut_1285_out;
            end
        end
        
        assign out_data[1285] = lut_1285_ff;
    end
    else begin : no_ff_1285
        assign out_data[1285] = lut_1285_out;
    end
    endgenerate
    
    
    
    // LUT : 1286
    wire [63:0] lut_1286_table = 64'b0000000000000010000000000000000000000010000000110000001000000011;
    wire [5:0] lut_1286_select = {
                             in_data[283],
                             in_data[699],
                             in_data[533],
                             in_data[127],
                             in_data[769],
                             in_data[667]};
    
    wire lut_1286_out = lut_1286_table[lut_1286_select];
    
    generate
    if ( USE_REG ) begin : ff_1286
        reg   lut_1286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1286_ff <= lut_1286_out;
            end
        end
        
        assign out_data[1286] = lut_1286_ff;
    end
    else begin : no_ff_1286
        assign out_data[1286] = lut_1286_out;
    end
    endgenerate
    
    
    
    // LUT : 1287
    wire [63:0] lut_1287_table = 64'b0000111100001111000011110000111100001111000011110000111100001111;
    wire [5:0] lut_1287_select = {
                             in_data[393],
                             in_data[0],
                             in_data[51],
                             in_data[213],
                             in_data[297],
                             in_data[39]};
    
    wire lut_1287_out = lut_1287_table[lut_1287_select];
    
    generate
    if ( USE_REG ) begin : ff_1287
        reg   lut_1287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1287_ff <= lut_1287_out;
            end
        end
        
        assign out_data[1287] = lut_1287_ff;
    end
    else begin : no_ff_1287
        assign out_data[1287] = lut_1287_out;
    end
    endgenerate
    
    
    
    // LUT : 1288
    wire [63:0] lut_1288_table = 64'b1010101010101010111110101010101011111010101010101111111111111010;
    wire [5:0] lut_1288_select = {
                             in_data[643],
                             in_data[228],
                             in_data[709],
                             in_data[430],
                             in_data[585],
                             in_data[427]};
    
    wire lut_1288_out = lut_1288_table[lut_1288_select];
    
    generate
    if ( USE_REG ) begin : ff_1288
        reg   lut_1288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1288_ff <= lut_1288_out;
            end
        end
        
        assign out_data[1288] = lut_1288_ff;
    end
    else begin : no_ff_1288
        assign out_data[1288] = lut_1288_out;
    end
    endgenerate
    
    
    
    // LUT : 1289
    wire [63:0] lut_1289_table = 64'b0000001100000011000011110000111100000011000000010000111100001111;
    wire [5:0] lut_1289_select = {
                             in_data[30],
                             in_data[631],
                             in_data[198],
                             in_data[149],
                             in_data[295],
                             in_data[449]};
    
    wire lut_1289_out = lut_1289_table[lut_1289_select];
    
    generate
    if ( USE_REG ) begin : ff_1289
        reg   lut_1289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1289_ff <= lut_1289_out;
            end
        end
        
        assign out_data[1289] = lut_1289_ff;
    end
    else begin : no_ff_1289
        assign out_data[1289] = lut_1289_out;
    end
    endgenerate
    
    
    
    // LUT : 1290
    wire [63:0] lut_1290_table = 64'b0000010100000101000001010000010100000101000001010000010100000101;
    wire [5:0] lut_1290_select = {
                             in_data[222],
                             in_data[109],
                             in_data[729],
                             in_data[227],
                             in_data[29],
                             in_data[597]};
    
    wire lut_1290_out = lut_1290_table[lut_1290_select];
    
    generate
    if ( USE_REG ) begin : ff_1290
        reg   lut_1290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1290_ff <= lut_1290_out;
            end
        end
        
        assign out_data[1290] = lut_1290_ff;
    end
    else begin : no_ff_1290
        assign out_data[1290] = lut_1290_out;
    end
    endgenerate
    
    
    
    // LUT : 1291
    wire [63:0] lut_1291_table = 64'b0000000000000000000001010000010100000101000001010101111100000101;
    wire [5:0] lut_1291_select = {
                             in_data[194],
                             in_data[221],
                             in_data[395],
                             in_data[555],
                             in_data[11],
                             in_data[578]};
    
    wire lut_1291_out = lut_1291_table[lut_1291_select];
    
    generate
    if ( USE_REG ) begin : ff_1291
        reg   lut_1291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1291_ff <= lut_1291_out;
            end
        end
        
        assign out_data[1291] = lut_1291_ff;
    end
    else begin : no_ff_1291
        assign out_data[1291] = lut_1291_out;
    end
    endgenerate
    
    
    
    // LUT : 1292
    wire [63:0] lut_1292_table = 64'b1111111111111101111111111111110111111101010101001111110101010100;
    wire [5:0] lut_1292_select = {
                             in_data[249],
                             in_data[35],
                             in_data[360],
                             in_data[245],
                             in_data[556],
                             in_data[664]};
    
    wire lut_1292_out = lut_1292_table[lut_1292_select];
    
    generate
    if ( USE_REG ) begin : ff_1292
        reg   lut_1292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1292_ff <= lut_1292_out;
            end
        end
        
        assign out_data[1292] = lut_1292_ff;
    end
    else begin : no_ff_1292
        assign out_data[1292] = lut_1292_out;
    end
    endgenerate
    
    
    
    // LUT : 1293
    wire [63:0] lut_1293_table = 64'b1110111111111111111011111111111100001100000011000000110000001100;
    wire [5:0] lut_1293_select = {
                             in_data[433],
                             in_data[615],
                             in_data[642],
                             in_data[527],
                             in_data[269],
                             in_data[735]};
    
    wire lut_1293_out = lut_1293_table[lut_1293_select];
    
    generate
    if ( USE_REG ) begin : ff_1293
        reg   lut_1293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1293_ff <= lut_1293_out;
            end
        end
        
        assign out_data[1293] = lut_1293_ff;
    end
    else begin : no_ff_1293
        assign out_data[1293] = lut_1293_out;
    end
    endgenerate
    
    
    
    // LUT : 1294
    wire [63:0] lut_1294_table = 64'b0000000000000000000011110010011100000000000000001010111110101111;
    wire [5:0] lut_1294_select = {
                             in_data[410],
                             in_data[469],
                             in_data[117],
                             in_data[529],
                             in_data[24],
                             in_data[381]};
    
    wire lut_1294_out = lut_1294_table[lut_1294_select];
    
    generate
    if ( USE_REG ) begin : ff_1294
        reg   lut_1294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1294_ff <= lut_1294_out;
            end
        end
        
        assign out_data[1294] = lut_1294_ff;
    end
    else begin : no_ff_1294
        assign out_data[1294] = lut_1294_out;
    end
    endgenerate
    
    
    
    // LUT : 1295
    wire [63:0] lut_1295_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1295_select = {
                             in_data[629],
                             in_data[418],
                             in_data[441],
                             in_data[738],
                             in_data[296],
                             in_data[516]};
    
    wire lut_1295_out = lut_1295_table[lut_1295_select];
    
    generate
    if ( USE_REG ) begin : ff_1295
        reg   lut_1295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1295_ff <= lut_1295_out;
            end
        end
        
        assign out_data[1295] = lut_1295_ff;
    end
    else begin : no_ff_1295
        assign out_data[1295] = lut_1295_out;
    end
    endgenerate
    
    
    
    // LUT : 1296
    wire [63:0] lut_1296_table = 64'b0000001100110011000000010001001100001011001100110000101100010011;
    wire [5:0] lut_1296_select = {
                             in_data[105],
                             in_data[111],
                             in_data[547],
                             in_data[128],
                             in_data[292],
                             in_data[359]};
    
    wire lut_1296_out = lut_1296_table[lut_1296_select];
    
    generate
    if ( USE_REG ) begin : ff_1296
        reg   lut_1296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1296_ff <= lut_1296_out;
            end
        end
        
        assign out_data[1296] = lut_1296_ff;
    end
    else begin : no_ff_1296
        assign out_data[1296] = lut_1296_out;
    end
    endgenerate
    
    
    
    // LUT : 1297
    wire [63:0] lut_1297_table = 64'b0011001011101000001100111110111011110011111111101111001111111111;
    wire [5:0] lut_1297_select = {
                             in_data[375],
                             in_data[50],
                             in_data[298],
                             in_data[665],
                             in_data[302],
                             in_data[123]};
    
    wire lut_1297_out = lut_1297_table[lut_1297_select];
    
    generate
    if ( USE_REG ) begin : ff_1297
        reg   lut_1297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1297_ff <= lut_1297_out;
            end
        end
        
        assign out_data[1297] = lut_1297_ff;
    end
    else begin : no_ff_1297
        assign out_data[1297] = lut_1297_out;
    end
    endgenerate
    
    
    
    // LUT : 1298
    wire [63:0] lut_1298_table = 64'b0100010011001100111111111111111101001100010011001111111111111111;
    wire [5:0] lut_1298_select = {
                             in_data[646],
                             in_data[356],
                             in_data[741],
                             in_data[133],
                             in_data[285],
                             in_data[568]};
    
    wire lut_1298_out = lut_1298_table[lut_1298_select];
    
    generate
    if ( USE_REG ) begin : ff_1298
        reg   lut_1298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1298_ff <= lut_1298_out;
            end
        end
        
        assign out_data[1298] = lut_1298_ff;
    end
    else begin : no_ff_1298
        assign out_data[1298] = lut_1298_out;
    end
    endgenerate
    
    
    
    // LUT : 1299
    wire [63:0] lut_1299_table = 64'b1010101001011010111110101111000010101010010110101111101011111010;
    wire [5:0] lut_1299_select = {
                             in_data[18],
                             in_data[549],
                             in_data[160],
                             in_data[436],
                             in_data[698],
                             in_data[272]};
    
    wire lut_1299_out = lut_1299_table[lut_1299_select];
    
    generate
    if ( USE_REG ) begin : ff_1299
        reg   lut_1299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1299_ff <= lut_1299_out;
            end
        end
        
        assign out_data[1299] = lut_1299_ff;
    end
    else begin : no_ff_1299
        assign out_data[1299] = lut_1299_out;
    end
    endgenerate
    
    
    
    // LUT : 1300
    wire [63:0] lut_1300_table = 64'b1111111111110000111111111111000011111111111100001111111111110000;
    wire [5:0] lut_1300_select = {
                             in_data[307],
                             in_data[448],
                             in_data[746],
                             in_data[237],
                             in_data[93],
                             in_data[780]};
    
    wire lut_1300_out = lut_1300_table[lut_1300_select];
    
    generate
    if ( USE_REG ) begin : ff_1300
        reg   lut_1300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1300_ff <= lut_1300_out;
            end
        end
        
        assign out_data[1300] = lut_1300_ff;
    end
    else begin : no_ff_1300
        assign out_data[1300] = lut_1300_out;
    end
    endgenerate
    
    
    
    // LUT : 1301
    wire [63:0] lut_1301_table = 64'b1101111111011111110011011100110111111111110111111100110001001100;
    wire [5:0] lut_1301_select = {
                             in_data[775],
                             in_data[507],
                             in_data[223],
                             in_data[424],
                             in_data[123],
                             in_data[687]};
    
    wire lut_1301_out = lut_1301_table[lut_1301_select];
    
    generate
    if ( USE_REG ) begin : ff_1301
        reg   lut_1301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1301_ff <= lut_1301_out;
            end
        end
        
        assign out_data[1301] = lut_1301_ff;
    end
    else begin : no_ff_1301
        assign out_data[1301] = lut_1301_out;
    end
    endgenerate
    
    
    
    // LUT : 1302
    wire [63:0] lut_1302_table = 64'b1111111101110111111111110101010111111111011101111111111101010101;
    wire [5:0] lut_1302_select = {
                             in_data[645],
                             in_data[471],
                             in_data[554],
                             in_data[506],
                             in_data[721],
                             in_data[268]};
    
    wire lut_1302_out = lut_1302_table[lut_1302_select];
    
    generate
    if ( USE_REG ) begin : ff_1302
        reg   lut_1302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1302_ff <= lut_1302_out;
            end
        end
        
        assign out_data[1302] = lut_1302_ff;
    end
    else begin : no_ff_1302
        assign out_data[1302] = lut_1302_out;
    end
    endgenerate
    
    
    
    // LUT : 1303
    wire [63:0] lut_1303_table = 64'b1111111100100010111111110010001011111111101010101111111110101010;
    wire [5:0] lut_1303_select = {
                             in_data[354],
                             in_data[144],
                             in_data[387],
                             in_data[54],
                             in_data[743],
                             in_data[410]};
    
    wire lut_1303_out = lut_1303_table[lut_1303_select];
    
    generate
    if ( USE_REG ) begin : ff_1303
        reg   lut_1303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1303_ff <= lut_1303_out;
            end
        end
        
        assign out_data[1303] = lut_1303_ff;
    end
    else begin : no_ff_1303
        assign out_data[1303] = lut_1303_out;
    end
    endgenerate
    
    
    
    // LUT : 1304
    wire [63:0] lut_1304_table = 64'b0000000011111111000000001111111100000000110111010100110011111111;
    wire [5:0] lut_1304_select = {
                             in_data[516],
                             in_data[484],
                             in_data[626],
                             in_data[25],
                             in_data[389],
                             in_data[13]};
    
    wire lut_1304_out = lut_1304_table[lut_1304_select];
    
    generate
    if ( USE_REG ) begin : ff_1304
        reg   lut_1304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1304_ff <= lut_1304_out;
            end
        end
        
        assign out_data[1304] = lut_1304_ff;
    end
    else begin : no_ff_1304
        assign out_data[1304] = lut_1304_out;
    end
    endgenerate
    
    
    
    // LUT : 1305
    wire [63:0] lut_1305_table = 64'b1111111100110011011101110010001111111111001100110111011100110011;
    wire [5:0] lut_1305_select = {
                             in_data[167],
                             in_data[479],
                             in_data[480],
                             in_data[42],
                             in_data[398],
                             in_data[269]};
    
    wire lut_1305_out = lut_1305_table[lut_1305_select];
    
    generate
    if ( USE_REG ) begin : ff_1305
        reg   lut_1305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1305_ff <= lut_1305_out;
            end
        end
        
        assign out_data[1305] = lut_1305_ff;
    end
    else begin : no_ff_1305
        assign out_data[1305] = lut_1305_out;
    end
    endgenerate
    
    
    
    // LUT : 1306
    wire [63:0] lut_1306_table = 64'b1101010111010000111101011101000111111101111101011111110111110101;
    wire [5:0] lut_1306_select = {
                             in_data[218],
                             in_data[765],
                             in_data[106],
                             in_data[100],
                             in_data[403],
                             in_data[628]};
    
    wire lut_1306_out = lut_1306_table[lut_1306_select];
    
    generate
    if ( USE_REG ) begin : ff_1306
        reg   lut_1306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1306_ff <= lut_1306_out;
            end
        end
        
        assign out_data[1306] = lut_1306_ff;
    end
    else begin : no_ff_1306
        assign out_data[1306] = lut_1306_out;
    end
    endgenerate
    
    
    
    // LUT : 1307
    wire [63:0] lut_1307_table = 64'b0101011100010101000000000000000001010101010101010000000000000001;
    wire [5:0] lut_1307_select = {
                             in_data[615],
                             in_data[740],
                             in_data[753],
                             in_data[48],
                             in_data[612],
                             in_data[564]};
    
    wire lut_1307_out = lut_1307_table[lut_1307_select];
    
    generate
    if ( USE_REG ) begin : ff_1307
        reg   lut_1307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1307_ff <= lut_1307_out;
            end
        end
        
        assign out_data[1307] = lut_1307_ff;
    end
    else begin : no_ff_1307
        assign out_data[1307] = lut_1307_out;
    end
    endgenerate
    
    
    
    // LUT : 1308
    wire [63:0] lut_1308_table = 64'b1000000010000000000000000000000000000001000000000000001100000000;
    wire [5:0] lut_1308_select = {
                             in_data[663],
                             in_data[146],
                             in_data[375],
                             in_data[660],
                             in_data[287],
                             in_data[386]};
    
    wire lut_1308_out = lut_1308_table[lut_1308_select];
    
    generate
    if ( USE_REG ) begin : ff_1308
        reg   lut_1308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1308_ff <= lut_1308_out;
            end
        end
        
        assign out_data[1308] = lut_1308_ff;
    end
    else begin : no_ff_1308
        assign out_data[1308] = lut_1308_out;
    end
    endgenerate
    
    
    
    // LUT : 1309
    wire [63:0] lut_1309_table = 64'b1111111101010101110111110101010100000000010101010000000001010101;
    wire [5:0] lut_1309_select = {
                             in_data[383],
                             in_data[168],
                             in_data[517],
                             in_data[773],
                             in_data[111],
                             in_data[605]};
    
    wire lut_1309_out = lut_1309_table[lut_1309_select];
    
    generate
    if ( USE_REG ) begin : ff_1309
        reg   lut_1309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1309_ff <= lut_1309_out;
            end
        end
        
        assign out_data[1309] = lut_1309_ff;
    end
    else begin : no_ff_1309
        assign out_data[1309] = lut_1309_out;
    end
    endgenerate
    
    
    
    // LUT : 1310
    wire [63:0] lut_1310_table = 64'b1100111111001111111011111110111100001100000011000000110000001100;
    wire [5:0] lut_1310_select = {
                             in_data[600],
                             in_data[150],
                             in_data[722],
                             in_data[492],
                             in_data[667],
                             in_data[716]};
    
    wire lut_1310_out = lut_1310_table[lut_1310_select];
    
    generate
    if ( USE_REG ) begin : ff_1310
        reg   lut_1310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1310_ff <= lut_1310_out;
            end
        end
        
        assign out_data[1310] = lut_1310_ff;
    end
    else begin : no_ff_1310
        assign out_data[1310] = lut_1310_out;
    end
    endgenerate
    
    
    
    // LUT : 1311
    wire [63:0] lut_1311_table = 64'b0000001100000011000011110000011100110000000100000011001100110011;
    wire [5:0] lut_1311_select = {
                             in_data[158],
                             in_data[341],
                             in_data[197],
                             in_data[601],
                             in_data[510],
                             in_data[676]};
    
    wire lut_1311_out = lut_1311_table[lut_1311_select];
    
    generate
    if ( USE_REG ) begin : ff_1311
        reg   lut_1311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1311_ff <= lut_1311_out;
            end
        end
        
        assign out_data[1311] = lut_1311_ff;
    end
    else begin : no_ff_1311
        assign out_data[1311] = lut_1311_out;
    end
    endgenerate
    
    
    
    // LUT : 1312
    wire [63:0] lut_1312_table = 64'b0000000000000000000000000000000000000000000000000101010101010101;
    wire [5:0] lut_1312_select = {
                             in_data[388],
                             in_data[414],
                             in_data[732],
                             in_data[557],
                             in_data[89],
                             in_data[467]};
    
    wire lut_1312_out = lut_1312_table[lut_1312_select];
    
    generate
    if ( USE_REG ) begin : ff_1312
        reg   lut_1312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1312_ff <= lut_1312_out;
            end
        end
        
        assign out_data[1312] = lut_1312_ff;
    end
    else begin : no_ff_1312
        assign out_data[1312] = lut_1312_out;
    end
    endgenerate
    
    
    
    // LUT : 1313
    wire [63:0] lut_1313_table = 64'b1111111111111111101010111111111110101010101010111010000010100010;
    wire [5:0] lut_1313_select = {
                             in_data[219],
                             in_data[686],
                             in_data[343],
                             in_data[549],
                             in_data[254],
                             in_data[207]};
    
    wire lut_1313_out = lut_1313_table[lut_1313_select];
    
    generate
    if ( USE_REG ) begin : ff_1313
        reg   lut_1313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1313_ff <= lut_1313_out;
            end
        end
        
        assign out_data[1313] = lut_1313_ff;
    end
    else begin : no_ff_1313
        assign out_data[1313] = lut_1313_out;
    end
    endgenerate
    
    
    
    // LUT : 1314
    wire [63:0] lut_1314_table = 64'b1000100010001100100010011000110110001101100011001000110110001100;
    wire [5:0] lut_1314_select = {
                             in_data[573],
                             in_data[113],
                             in_data[101],
                             in_data[267],
                             in_data[515],
                             in_data[460]};
    
    wire lut_1314_out = lut_1314_table[lut_1314_select];
    
    generate
    if ( USE_REG ) begin : ff_1314
        reg   lut_1314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1314_ff <= lut_1314_out;
            end
        end
        
        assign out_data[1314] = lut_1314_ff;
    end
    else begin : no_ff_1314
        assign out_data[1314] = lut_1314_out;
    end
    endgenerate
    
    
    
    // LUT : 1315
    wire [63:0] lut_1315_table = 64'b0000000000000000111100101110001100000000000000000000001111001111;
    wire [5:0] lut_1315_select = {
                             in_data[332],
                             in_data[322],
                             in_data[171],
                             in_data[160],
                             in_data[103],
                             in_data[252]};
    
    wire lut_1315_out = lut_1315_table[lut_1315_select];
    
    generate
    if ( USE_REG ) begin : ff_1315
        reg   lut_1315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1315_ff <= lut_1315_out;
            end
        end
        
        assign out_data[1315] = lut_1315_ff;
    end
    else begin : no_ff_1315
        assign out_data[1315] = lut_1315_out;
    end
    endgenerate
    
    
    
    // LUT : 1316
    wire [63:0] lut_1316_table = 64'b1111111111111111110011001100110111111111111111110000000000000000;
    wire [5:0] lut_1316_select = {
                             in_data[125],
                             in_data[294],
                             in_data[726],
                             in_data[280],
                             in_data[352],
                             in_data[82]};
    
    wire lut_1316_out = lut_1316_table[lut_1316_select];
    
    generate
    if ( USE_REG ) begin : ff_1316
        reg   lut_1316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1316_ff <= lut_1316_out;
            end
        end
        
        assign out_data[1316] = lut_1316_ff;
    end
    else begin : no_ff_1316
        assign out_data[1316] = lut_1316_out;
    end
    endgenerate
    
    
    
    // LUT : 1317
    wire [63:0] lut_1317_table = 64'b1111111111110000111111111111000011111111111100001111111111110000;
    wire [5:0] lut_1317_select = {
                             in_data[342],
                             in_data[61],
                             in_data[579],
                             in_data[193],
                             in_data[199],
                             in_data[758]};
    
    wire lut_1317_out = lut_1317_table[lut_1317_select];
    
    generate
    if ( USE_REG ) begin : ff_1317
        reg   lut_1317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1317_ff <= lut_1317_out;
            end
        end
        
        assign out_data[1317] = lut_1317_ff;
    end
    else begin : no_ff_1317
        assign out_data[1317] = lut_1317_out;
    end
    endgenerate
    
    
    
    // LUT : 1318
    wire [63:0] lut_1318_table = 64'b1011111110111110101111111011111100001100010011000000010100000101;
    wire [5:0] lut_1318_select = {
                             in_data[303],
                             in_data[576],
                             in_data[723],
                             in_data[128],
                             in_data[372],
                             in_data[513]};
    
    wire lut_1318_out = lut_1318_table[lut_1318_select];
    
    generate
    if ( USE_REG ) begin : ff_1318
        reg   lut_1318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1318_ff <= lut_1318_out;
            end
        end
        
        assign out_data[1318] = lut_1318_ff;
    end
    else begin : no_ff_1318
        assign out_data[1318] = lut_1318_out;
    end
    endgenerate
    
    
    
    // LUT : 1319
    wire [63:0] lut_1319_table = 64'b0000000000000000000000000000000000010011000100010001000100010001;
    wire [5:0] lut_1319_select = {
                             in_data[245],
                             in_data[262],
                             in_data[32],
                             in_data[16],
                             in_data[261],
                             in_data[272]};
    
    wire lut_1319_out = lut_1319_table[lut_1319_select];
    
    generate
    if ( USE_REG ) begin : ff_1319
        reg   lut_1319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1319_ff <= lut_1319_out;
            end
        end
        
        assign out_data[1319] = lut_1319_ff;
    end
    else begin : no_ff_1319
        assign out_data[1319] = lut_1319_out;
    end
    endgenerate
    
    
    
    // LUT : 1320
    wire [63:0] lut_1320_table = 64'b1111000010100000111111111111010111110000101000001111111111110100;
    wire [5:0] lut_1320_select = {
                             in_data[19],
                             in_data[511],
                             in_data[119],
                             in_data[323],
                             in_data[35],
                             in_data[329]};
    
    wire lut_1320_out = lut_1320_table[lut_1320_select];
    
    generate
    if ( USE_REG ) begin : ff_1320
        reg   lut_1320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1320_ff <= lut_1320_out;
            end
        end
        
        assign out_data[1320] = lut_1320_ff;
    end
    else begin : no_ff_1320
        assign out_data[1320] = lut_1320_out;
    end
    endgenerate
    
    
    
    // LUT : 1321
    wire [63:0] lut_1321_table = 64'b0010111100101110001011110010111100101111101011110010111110001111;
    wire [5:0] lut_1321_select = {
                             in_data[115],
                             in_data[50],
                             in_data[501],
                             in_data[521],
                             in_data[529],
                             in_data[520]};
    
    wire lut_1321_out = lut_1321_table[lut_1321_select];
    
    generate
    if ( USE_REG ) begin : ff_1321
        reg   lut_1321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1321_ff <= lut_1321_out;
            end
        end
        
        assign out_data[1321] = lut_1321_ff;
    end
    else begin : no_ff_1321
        assign out_data[1321] = lut_1321_out;
    end
    endgenerate
    
    
    
    // LUT : 1322
    wire [63:0] lut_1322_table = 64'b0000000000000000000000000000000011010101110101011111101111111010;
    wire [5:0] lut_1322_select = {
                             in_data[592],
                             in_data[183],
                             in_data[56],
                             in_data[367],
                             in_data[99],
                             in_data[680]};
    
    wire lut_1322_out = lut_1322_table[lut_1322_select];
    
    generate
    if ( USE_REG ) begin : ff_1322
        reg   lut_1322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1322_ff <= lut_1322_out;
            end
        end
        
        assign out_data[1322] = lut_1322_ff;
    end
    else begin : no_ff_1322
        assign out_data[1322] = lut_1322_out;
    end
    endgenerate
    
    
    
    // LUT : 1323
    wire [63:0] lut_1323_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1323_select = {
                             in_data[700],
                             in_data[688],
                             in_data[558],
                             in_data[36],
                             in_data[324],
                             in_data[338]};
    
    wire lut_1323_out = lut_1323_table[lut_1323_select];
    
    generate
    if ( USE_REG ) begin : ff_1323
        reg   lut_1323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1323_ff <= lut_1323_out;
            end
        end
        
        assign out_data[1323] = lut_1323_ff;
    end
    else begin : no_ff_1323
        assign out_data[1323] = lut_1323_out;
    end
    endgenerate
    
    
    
    // LUT : 1324
    wire [63:0] lut_1324_table = 64'b0000000000000000000000000000000000000000111111111111111111111111;
    wire [5:0] lut_1324_select = {
                             in_data[401],
                             in_data[68],
                             in_data[487],
                             in_data[309],
                             in_data[79],
                             in_data[365]};
    
    wire lut_1324_out = lut_1324_table[lut_1324_select];
    
    generate
    if ( USE_REG ) begin : ff_1324
        reg   lut_1324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1324_ff <= lut_1324_out;
            end
        end
        
        assign out_data[1324] = lut_1324_ff;
    end
    else begin : no_ff_1324
        assign out_data[1324] = lut_1324_out;
    end
    endgenerate
    
    
    
    // LUT : 1325
    wire [63:0] lut_1325_table = 64'b0000001100000001000000000000000000000011000000010000000100010001;
    wire [5:0] lut_1325_select = {
                             in_data[710],
                             in_data[653],
                             in_data[96],
                             in_data[627],
                             in_data[148],
                             in_data[526]};
    
    wire lut_1325_out = lut_1325_table[lut_1325_select];
    
    generate
    if ( USE_REG ) begin : ff_1325
        reg   lut_1325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1325_ff <= lut_1325_out;
            end
        end
        
        assign out_data[1325] = lut_1325_ff;
    end
    else begin : no_ff_1325
        assign out_data[1325] = lut_1325_out;
    end
    endgenerate
    
    
    
    // LUT : 1326
    wire [63:0] lut_1326_table = 64'b0000111100001111000011110000111100001110000011100000111000001111;
    wire [5:0] lut_1326_select = {
                             in_data[143],
                             in_data[781],
                             in_data[90],
                             in_data[156],
                             in_data[531],
                             in_data[381]};
    
    wire lut_1326_out = lut_1326_table[lut_1326_select];
    
    generate
    if ( USE_REG ) begin : ff_1326
        reg   lut_1326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1326_ff <= lut_1326_out;
            end
        end
        
        assign out_data[1326] = lut_1326_ff;
    end
    else begin : no_ff_1326
        assign out_data[1326] = lut_1326_out;
    end
    endgenerate
    
    
    
    // LUT : 1327
    wire [63:0] lut_1327_table = 64'b1111111111111111111111111111111100000000000000001111111111111111;
    wire [5:0] lut_1327_select = {
                             in_data[425],
                             in_data[597],
                             in_data[105],
                             in_data[306],
                             in_data[310],
                             in_data[613]};
    
    wire lut_1327_out = lut_1327_table[lut_1327_select];
    
    generate
    if ( USE_REG ) begin : ff_1327
        reg   lut_1327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1327_ff <= lut_1327_out;
            end
        end
        
        assign out_data[1327] = lut_1327_ff;
    end
    else begin : no_ff_1327
        assign out_data[1327] = lut_1327_out;
    end
    endgenerate
    
    
    
    // LUT : 1328
    wire [63:0] lut_1328_table = 64'b0000000001010000000000000101000001010000010101010101000001010101;
    wire [5:0] lut_1328_select = {
                             in_data[351],
                             in_data[20],
                             in_data[611],
                             in_data[69],
                             in_data[226],
                             in_data[555]};
    
    wire lut_1328_out = lut_1328_table[lut_1328_select];
    
    generate
    if ( USE_REG ) begin : ff_1328
        reg   lut_1328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1328_ff <= lut_1328_out;
            end
        end
        
        assign out_data[1328] = lut_1328_ff;
    end
    else begin : no_ff_1328
        assign out_data[1328] = lut_1328_out;
    end
    endgenerate
    
    
    
    // LUT : 1329
    wire [63:0] lut_1329_table = 64'b0101010101010101010101010101010101010101010101010101010101010101;
    wire [5:0] lut_1329_select = {
                             in_data[704],
                             in_data[46],
                             in_data[675],
                             in_data[629],
                             in_data[644],
                             in_data[177]};
    
    wire lut_1329_out = lut_1329_table[lut_1329_select];
    
    generate
    if ( USE_REG ) begin : ff_1329
        reg   lut_1329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1329_ff <= lut_1329_out;
            end
        end
        
        assign out_data[1329] = lut_1329_ff;
    end
    else begin : no_ff_1329
        assign out_data[1329] = lut_1329_out;
    end
    endgenerate
    
    
    
    // LUT : 1330
    wire [63:0] lut_1330_table = 64'b0000010100001000000001010000000011111111100011100101111100001000;
    wire [5:0] lut_1330_select = {
                             in_data[621],
                             in_data[78],
                             in_data[458],
                             in_data[735],
                             in_data[138],
                             in_data[134]};
    
    wire lut_1330_out = lut_1330_table[lut_1330_select];
    
    generate
    if ( USE_REG ) begin : ff_1330
        reg   lut_1330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1330_ff <= lut_1330_out;
            end
        end
        
        assign out_data[1330] = lut_1330_ff;
    end
    else begin : no_ff_1330
        assign out_data[1330] = lut_1330_out;
    end
    endgenerate
    
    
    
    // LUT : 1331
    wire [63:0] lut_1331_table = 64'b1111111111111111111110001111100011111111111111111111100011110000;
    wire [5:0] lut_1331_select = {
                             in_data[783],
                             in_data[413],
                             in_data[444],
                             in_data[244],
                             in_data[209],
                             in_data[649]};
    
    wire lut_1331_out = lut_1331_table[lut_1331_select];
    
    generate
    if ( USE_REG ) begin : ff_1331
        reg   lut_1331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1331_ff <= lut_1331_out;
            end
        end
        
        assign out_data[1331] = lut_1331_ff;
    end
    else begin : no_ff_1331
        assign out_data[1331] = lut_1331_out;
    end
    endgenerate
    
    
    
    // LUT : 1332
    wire [63:0] lut_1332_table = 64'b1111111100001111111111110000111111111111000011101111111100001110;
    wire [5:0] lut_1332_select = {
                             in_data[563],
                             in_data[561],
                             in_data[464],
                             in_data[263],
                             in_data[356],
                             in_data[145]};
    
    wire lut_1332_out = lut_1332_table[lut_1332_select];
    
    generate
    if ( USE_REG ) begin : ff_1332
        reg   lut_1332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1332_ff <= lut_1332_out;
            end
        end
        
        assign out_data[1332] = lut_1332_ff;
    end
    else begin : no_ff_1332
        assign out_data[1332] = lut_1332_out;
    end
    endgenerate
    
    
    
    // LUT : 1333
    wire [63:0] lut_1333_table = 64'b0000000000000000000000000000000000001100000011000000111100001111;
    wire [5:0] lut_1333_select = {
                             in_data[607],
                             in_data[538],
                             in_data[586],
                             in_data[133],
                             in_data[584],
                             in_data[73]};
    
    wire lut_1333_out = lut_1333_table[lut_1333_select];
    
    generate
    if ( USE_REG ) begin : ff_1333
        reg   lut_1333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1333_ff <= lut_1333_out;
            end
        end
        
        assign out_data[1333] = lut_1333_ff;
    end
    else begin : no_ff_1333
        assign out_data[1333] = lut_1333_out;
    end
    endgenerate
    
    
    
    // LUT : 1334
    wire [63:0] lut_1334_table = 64'b1100111111111111111111111111111100001100000011000000110000001100;
    wire [5:0] lut_1334_select = {
                             in_data[357],
                             in_data[706],
                             in_data[598],
                             in_data[178],
                             in_data[313],
                             in_data[59]};
    
    wire lut_1334_out = lut_1334_table[lut_1334_select];
    
    generate
    if ( USE_REG ) begin : ff_1334
        reg   lut_1334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1334_ff <= lut_1334_out;
            end
        end
        
        assign out_data[1334] = lut_1334_ff;
    end
    else begin : no_ff_1334
        assign out_data[1334] = lut_1334_out;
    end
    endgenerate
    
    
    
    // LUT : 1335
    wire [63:0] lut_1335_table = 64'b1100111011001111010001000100010000110011001100110000000000000000;
    wire [5:0] lut_1335_select = {
                             in_data[259],
                             in_data[318],
                             in_data[198],
                             in_data[734],
                             in_data[638],
                             in_data[543]};
    
    wire lut_1335_out = lut_1335_table[lut_1335_select];
    
    generate
    if ( USE_REG ) begin : ff_1335
        reg   lut_1335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1335_ff <= lut_1335_out;
            end
        end
        
        assign out_data[1335] = lut_1335_ff;
    end
    else begin : no_ff_1335
        assign out_data[1335] = lut_1335_out;
    end
    endgenerate
    
    
    
    // LUT : 1336
    wire [63:0] lut_1336_table = 64'b0111111101110111011101110111011100010001000100010001000100010001;
    wire [5:0] lut_1336_select = {
                             in_data[684],
                             in_data[720],
                             in_data[222],
                             in_data[165],
                             in_data[498],
                             in_data[689]};
    
    wire lut_1336_out = lut_1336_table[lut_1336_select];
    
    generate
    if ( USE_REG ) begin : ff_1336
        reg   lut_1336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1336_ff <= lut_1336_out;
            end
        end
        
        assign out_data[1336] = lut_1336_ff;
    end
    else begin : no_ff_1336
        assign out_data[1336] = lut_1336_out;
    end
    endgenerate
    
    
    
    // LUT : 1337
    wire [63:0] lut_1337_table = 64'b0011001100000001001100110000000000110011000000110011001100000000;
    wire [5:0] lut_1337_select = {
                             in_data[763],
                             in_data[572],
                             in_data[320],
                             in_data[537],
                             in_data[124],
                             in_data[624]};
    
    wire lut_1337_out = lut_1337_table[lut_1337_select];
    
    generate
    if ( USE_REG ) begin : ff_1337
        reg   lut_1337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1337_ff <= lut_1337_out;
            end
        end
        
        assign out_data[1337] = lut_1337_ff;
    end
    else begin : no_ff_1337
        assign out_data[1337] = lut_1337_out;
    end
    endgenerate
    
    
    
    // LUT : 1338
    wire [63:0] lut_1338_table = 64'b1111111111111111111111111010111111111111101011111110111110001100;
    wire [5:0] lut_1338_select = {
                             in_data[714],
                             in_data[238],
                             in_data[249],
                             in_data[147],
                             in_data[312],
                             in_data[260]};
    
    wire lut_1338_out = lut_1338_table[lut_1338_select];
    
    generate
    if ( USE_REG ) begin : ff_1338
        reg   lut_1338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1338_ff <= lut_1338_out;
            end
        end
        
        assign out_data[1338] = lut_1338_ff;
    end
    else begin : no_ff_1338
        assign out_data[1338] = lut_1338_out;
    end
    endgenerate
    
    
    
    // LUT : 1339
    wire [63:0] lut_1339_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_1339_select = {
                             in_data[760],
                             in_data[437],
                             in_data[514],
                             in_data[83],
                             in_data[131],
                             in_data[392]};
    
    wire lut_1339_out = lut_1339_table[lut_1339_select];
    
    generate
    if ( USE_REG ) begin : ff_1339
        reg   lut_1339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1339_ff <= lut_1339_out;
            end
        end
        
        assign out_data[1339] = lut_1339_ff;
    end
    else begin : no_ff_1339
        assign out_data[1339] = lut_1339_out;
    end
    endgenerate
    
    
    
    // LUT : 1340
    wire [63:0] lut_1340_table = 64'b1010101010101010101010101010101011111111111111111111111111111111;
    wire [5:0] lut_1340_select = {
                             in_data[512],
                             in_data[637],
                             in_data[643],
                             in_data[552],
                             in_data[768],
                             in_data[192]};
    
    wire lut_1340_out = lut_1340_table[lut_1340_select];
    
    generate
    if ( USE_REG ) begin : ff_1340
        reg   lut_1340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1340_ff <= lut_1340_out;
            end
        end
        
        assign out_data[1340] = lut_1340_ff;
    end
    else begin : no_ff_1340
        assign out_data[1340] = lut_1340_out;
    end
    endgenerate
    
    
    
    // LUT : 1341
    wire [63:0] lut_1341_table = 64'b1111111111111111101010101000101011111111111111111010111010101010;
    wire [5:0] lut_1341_select = {
                             in_data[293],
                             in_data[407],
                             in_data[37],
                             in_data[200],
                             in_data[450],
                             in_data[678]};
    
    wire lut_1341_out = lut_1341_table[lut_1341_select];
    
    generate
    if ( USE_REG ) begin : ff_1341
        reg   lut_1341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1341_ff <= lut_1341_out;
            end
        end
        
        assign out_data[1341] = lut_1341_ff;
    end
    else begin : no_ff_1341
        assign out_data[1341] = lut_1341_out;
    end
    endgenerate
    
    
    
    // LUT : 1342
    wire [63:0] lut_1342_table = 64'b0000000000100010111111111111111100000000000000001010101010111011;
    wire [5:0] lut_1342_select = {
                             in_data[548],
                             in_data[379],
                             in_data[500],
                             in_data[142],
                             in_data[705],
                             in_data[652]};
    
    wire lut_1342_out = lut_1342_table[lut_1342_select];
    
    generate
    if ( USE_REG ) begin : ff_1342
        reg   lut_1342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1342_ff <= lut_1342_out;
            end
        end
        
        assign out_data[1342] = lut_1342_ff;
    end
    else begin : no_ff_1342
        assign out_data[1342] = lut_1342_out;
    end
    endgenerate
    
    
    
    // LUT : 1343
    wire [63:0] lut_1343_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1343_select = {
                             in_data[568],
                             in_data[540],
                             in_data[139],
                             in_data[185],
                             in_data[374],
                             in_data[583]};
    
    wire lut_1343_out = lut_1343_table[lut_1343_select];
    
    generate
    if ( USE_REG ) begin : ff_1343
        reg   lut_1343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1343_ff <= lut_1343_out;
            end
        end
        
        assign out_data[1343] = lut_1343_ff;
    end
    else begin : no_ff_1343
        assign out_data[1343] = lut_1343_out;
    end
    endgenerate
    
    
    
    // LUT : 1344
    wire [63:0] lut_1344_table = 64'b1111111111101101111111111110110111111111111011011111111111101101;
    wire [5:0] lut_1344_select = {
                             in_data[86],
                             in_data[761],
                             in_data[120],
                             in_data[608],
                             in_data[164],
                             in_data[292]};
    
    wire lut_1344_out = lut_1344_table[lut_1344_select];
    
    generate
    if ( USE_REG ) begin : ff_1344
        reg   lut_1344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1344_ff <= lut_1344_out;
            end
        end
        
        assign out_data[1344] = lut_1344_ff;
    end
    else begin : no_ff_1344
        assign out_data[1344] = lut_1344_out;
    end
    endgenerate
    
    
    
    // LUT : 1345
    wire [63:0] lut_1345_table = 64'b0000000000000000000000000000001100000000000000110000000000111111;
    wire [5:0] lut_1345_select = {
                             in_data[399],
                             in_data[75],
                             in_data[455],
                             in_data[416],
                             in_data[715],
                             in_data[141]};
    
    wire lut_1345_out = lut_1345_table[lut_1345_select];
    
    generate
    if ( USE_REG ) begin : ff_1345
        reg   lut_1345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1345_ff <= lut_1345_out;
            end
        end
        
        assign out_data[1345] = lut_1345_ff;
    end
    else begin : no_ff_1345
        assign out_data[1345] = lut_1345_out;
    end
    endgenerate
    
    
    
    // LUT : 1346
    wire [63:0] lut_1346_table = 64'b0000000000000000001000101011101100000000000000001111111111111111;
    wire [5:0] lut_1346_select = {
                             in_data[625],
                             in_data[349],
                             in_data[685],
                             in_data[212],
                             in_data[508],
                             in_data[229]};
    
    wire lut_1346_out = lut_1346_table[lut_1346_select];
    
    generate
    if ( USE_REG ) begin : ff_1346
        reg   lut_1346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1346_ff <= lut_1346_out;
            end
        end
        
        assign out_data[1346] = lut_1346_ff;
    end
    else begin : no_ff_1346
        assign out_data[1346] = lut_1346_out;
    end
    endgenerate
    
    
    
    // LUT : 1347
    wire [63:0] lut_1347_table = 64'b1111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_1347_select = {
                             in_data[250],
                             in_data[777],
                             in_data[92],
                             in_data[599],
                             in_data[683],
                             in_data[729]};
    
    wire lut_1347_out = lut_1347_table[lut_1347_select];
    
    generate
    if ( USE_REG ) begin : ff_1347
        reg   lut_1347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1347_ff <= lut_1347_out;
            end
        end
        
        assign out_data[1347] = lut_1347_ff;
    end
    else begin : no_ff_1347
        assign out_data[1347] = lut_1347_out;
    end
    endgenerate
    
    
    
    // LUT : 1348
    wire [63:0] lut_1348_table = 64'b0000000000000000000000001111111100000000000000000000000011111111;
    wire [5:0] lut_1348_select = {
                             in_data[362],
                             in_data[384],
                             in_data[553],
                             in_data[308],
                             in_data[196],
                             in_data[646]};
    
    wire lut_1348_out = lut_1348_table[lut_1348_select];
    
    generate
    if ( USE_REG ) begin : ff_1348
        reg   lut_1348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1348_ff <= lut_1348_out;
            end
        end
        
        assign out_data[1348] = lut_1348_ff;
    end
    else begin : no_ff_1348
        assign out_data[1348] = lut_1348_out;
    end
    endgenerate
    
    
    
    // LUT : 1349
    wire [63:0] lut_1349_table = 64'b0101110100000000110111010000110101010101000000000101010100001100;
    wire [5:0] lut_1349_select = {
                             in_data[641],
                             in_data[182],
                             in_data[355],
                             in_data[98],
                             in_data[570],
                             in_data[214]};
    
    wire lut_1349_out = lut_1349_table[lut_1349_select];
    
    generate
    if ( USE_REG ) begin : ff_1349
        reg   lut_1349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1349_ff <= lut_1349_out;
            end
        end
        
        assign out_data[1349] = lut_1349_ff;
    end
    else begin : no_ff_1349
        assign out_data[1349] = lut_1349_out;
    end
    endgenerate
    
    
    
    // LUT : 1350
    wire [63:0] lut_1350_table = 64'b0000000011110111000000000000000001010101111111110101010111111111;
    wire [5:0] lut_1350_select = {
                             in_data[574],
                             in_data[136],
                             in_data[465],
                             in_data[81],
                             in_data[33],
                             in_data[284]};
    
    wire lut_1350_out = lut_1350_table[lut_1350_select];
    
    generate
    if ( USE_REG ) begin : ff_1350
        reg   lut_1350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1350_ff <= lut_1350_out;
            end
        end
        
        assign out_data[1350] = lut_1350_ff;
    end
    else begin : no_ff_1350
        assign out_data[1350] = lut_1350_out;
    end
    endgenerate
    
    
    
    // LUT : 1351
    wire [63:0] lut_1351_table = 64'b0000000000000000110111011100111000000000000000001101110111011101;
    wire [5:0] lut_1351_select = {
                             in_data[712],
                             in_data[152],
                             in_data[4],
                             in_data[672],
                             in_data[299],
                             in_data[562]};
    
    wire lut_1351_out = lut_1351_table[lut_1351_select];
    
    generate
    if ( USE_REG ) begin : ff_1351
        reg   lut_1351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1351_ff <= lut_1351_out;
            end
        end
        
        assign out_data[1351] = lut_1351_ff;
    end
    else begin : no_ff_1351
        assign out_data[1351] = lut_1351_out;
    end
    endgenerate
    
    
    
    // LUT : 1352
    wire [63:0] lut_1352_table = 64'b0000000001011111000000000101111000001010010011110000101000011111;
    wire [5:0] lut_1352_select = {
                             in_data[380],
                             in_data[116],
                             in_data[231],
                             in_data[129],
                             in_data[673],
                             in_data[211]};
    
    wire lut_1352_out = lut_1352_table[lut_1352_select];
    
    generate
    if ( USE_REG ) begin : ff_1352
        reg   lut_1352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1352_ff <= lut_1352_out;
            end
        end
        
        assign out_data[1352] = lut_1352_ff;
    end
    else begin : no_ff_1352
        assign out_data[1352] = lut_1352_out;
    end
    endgenerate
    
    
    
    // LUT : 1353
    wire [63:0] lut_1353_table = 64'b0000000000000000000000000000000000000000000100000001000100110001;
    wire [5:0] lut_1353_select = {
                             in_data[151],
                             in_data[71],
                             in_data[217],
                             in_data[210],
                             in_data[633],
                             in_data[72]};
    
    wire lut_1353_out = lut_1353_table[lut_1353_select];
    
    generate
    if ( USE_REG ) begin : ff_1353
        reg   lut_1353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1353_ff <= lut_1353_out;
            end
        end
        
        assign out_data[1353] = lut_1353_ff;
    end
    else begin : no_ff_1353
        assign out_data[1353] = lut_1353_out;
    end
    endgenerate
    
    
    
    // LUT : 1354
    wire [63:0] lut_1354_table = 64'b0001000001010101000000000101010100010000010101010000000001010101;
    wire [5:0] lut_1354_select = {
                             in_data[18],
                             in_data[85],
                             in_data[466],
                             in_data[474],
                             in_data[420],
                             in_data[639]};
    
    wire lut_1354_out = lut_1354_table[lut_1354_select];
    
    generate
    if ( USE_REG ) begin : ff_1354
        reg   lut_1354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1354_ff <= lut_1354_out;
            end
        end
        
        assign out_data[1354] = lut_1354_ff;
    end
    else begin : no_ff_1354
        assign out_data[1354] = lut_1354_out;
    end
    endgenerate
    
    
    
    // LUT : 1355
    wire [63:0] lut_1355_table = 64'b0000000000000000000000000000000100000000000000000000000100000001;
    wire [5:0] lut_1355_select = {
                             in_data[587],
                             in_data[443],
                             in_data[77],
                             in_data[719],
                             in_data[94],
                             in_data[28]};
    
    wire lut_1355_out = lut_1355_table[lut_1355_select];
    
    generate
    if ( USE_REG ) begin : ff_1355
        reg   lut_1355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1355_ff <= lut_1355_out;
            end
        end
        
        assign out_data[1355] = lut_1355_ff;
    end
    else begin : no_ff_1355
        assign out_data[1355] = lut_1355_out;
    end
    endgenerate
    
    
    
    // LUT : 1356
    wire [63:0] lut_1356_table = 64'b1010000011100000111111111111111100000000111100001111111111111111;
    wire [5:0] lut_1356_select = {
                             in_data[348],
                             in_data[427],
                             in_data[186],
                             in_data[176],
                             in_data[609],
                             in_data[65]};
    
    wire lut_1356_out = lut_1356_table[lut_1356_select];
    
    generate
    if ( USE_REG ) begin : ff_1356
        reg   lut_1356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1356_ff <= lut_1356_out;
            end
        end
        
        assign out_data[1356] = lut_1356_ff;
    end
    else begin : no_ff_1356
        assign out_data[1356] = lut_1356_out;
    end
    endgenerate
    
    
    
    // LUT : 1357
    wire [63:0] lut_1357_table = 64'b0001011100000000000000110010001000110011000000001010001010111010;
    wire [5:0] lut_1357_select = {
                             in_data[290],
                             in_data[661],
                             in_data[630],
                             in_data[302],
                             in_data[172],
                             in_data[541]};
    
    wire lut_1357_out = lut_1357_table[lut_1357_select];
    
    generate
    if ( USE_REG ) begin : ff_1357
        reg   lut_1357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1357_ff <= lut_1357_out;
            end
        end
        
        assign out_data[1357] = lut_1357_ff;
    end
    else begin : no_ff_1357
        assign out_data[1357] = lut_1357_out;
    end
    endgenerate
    
    
    
    // LUT : 1358
    wire [63:0] lut_1358_table = 64'b1111000011110000111111111111111111110000111100001111111111111111;
    wire [5:0] lut_1358_select = {
                             in_data[616],
                             in_data[485],
                             in_data[282],
                             in_data[189],
                             in_data[191],
                             in_data[642]};
    
    wire lut_1358_out = lut_1358_table[lut_1358_select];
    
    generate
    if ( USE_REG ) begin : ff_1358
        reg   lut_1358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1358_ff <= lut_1358_out;
            end
        end
        
        assign out_data[1358] = lut_1358_ff;
    end
    else begin : no_ff_1358
        assign out_data[1358] = lut_1358_out;
    end
    endgenerate
    
    
    
    // LUT : 1359
    wire [63:0] lut_1359_table = 64'b1111111111111111111111111111111111111100111111001111110011001100;
    wire [5:0] lut_1359_select = {
                             in_data[242],
                             in_data[556],
                             in_data[669],
                             in_data[640],
                             in_data[486],
                             in_data[109]};
    
    wire lut_1359_out = lut_1359_table[lut_1359_select];
    
    generate
    if ( USE_REG ) begin : ff_1359
        reg   lut_1359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1359_ff <= lut_1359_out;
            end
        end
        
        assign out_data[1359] = lut_1359_ff;
    end
    else begin : no_ff_1359
        assign out_data[1359] = lut_1359_out;
    end
    endgenerate
    
    
    
    // LUT : 1360
    wire [63:0] lut_1360_table = 64'b0000111100001111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_1360_select = {
                             in_data[662],
                             in_data[291],
                             in_data[80],
                             in_data[459],
                             in_data[449],
                             in_data[739]};
    
    wire lut_1360_out = lut_1360_table[lut_1360_select];
    
    generate
    if ( USE_REG ) begin : ff_1360
        reg   lut_1360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1360_ff <= lut_1360_out;
            end
        end
        
        assign out_data[1360] = lut_1360_ff;
    end
    else begin : no_ff_1360
        assign out_data[1360] = lut_1360_out;
    end
    endgenerate
    
    
    
    // LUT : 1361
    wire [63:0] lut_1361_table = 64'b1111101010100000111111111111111110100000100000001111101011111010;
    wire [5:0] lut_1361_select = {
                             in_data[206],
                             in_data[664],
                             in_data[40],
                             in_data[279],
                             in_data[762],
                             in_data[745]};
    
    wire lut_1361_out = lut_1361_table[lut_1361_select];
    
    generate
    if ( USE_REG ) begin : ff_1361
        reg   lut_1361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1361_ff <= lut_1361_out;
            end
        end
        
        assign out_data[1361] = lut_1361_ff;
    end
    else begin : no_ff_1361
        assign out_data[1361] = lut_1361_out;
    end
    endgenerate
    
    
    
    // LUT : 1362
    wire [63:0] lut_1362_table = 64'b1111010111111111000100001111010111110101111111110000000011110101;
    wire [5:0] lut_1362_select = {
                             in_data[84],
                             in_data[95],
                             in_data[273],
                             in_data[175],
                             in_data[49],
                             in_data[339]};
    
    wire lut_1362_out = lut_1362_table[lut_1362_select];
    
    generate
    if ( USE_REG ) begin : ff_1362
        reg   lut_1362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1362_ff <= lut_1362_out;
            end
        end
        
        assign out_data[1362] = lut_1362_ff;
    end
    else begin : no_ff_1362
        assign out_data[1362] = lut_1362_out;
    end
    endgenerate
    
    
    
    // LUT : 1363
    wire [63:0] lut_1363_table = 64'b0000000000000000000011110000111000000000000000000000111100001111;
    wire [5:0] lut_1363_select = {
                             in_data[224],
                             in_data[692],
                             in_data[536],
                             in_data[622],
                             in_data[0],
                             in_data[335]};
    
    wire lut_1363_out = lut_1363_table[lut_1363_select];
    
    generate
    if ( USE_REG ) begin : ff_1363
        reg   lut_1363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1363_ff <= lut_1363_out;
            end
        end
        
        assign out_data[1363] = lut_1363_ff;
    end
    else begin : no_ff_1363
        assign out_data[1363] = lut_1363_out;
    end
    endgenerate
    
    
    
    // LUT : 1364
    wire [63:0] lut_1364_table = 64'b1111111110101110111111111010101011111111101011101111111110101110;
    wire [5:0] lut_1364_select = {
                             in_data[772],
                             in_data[9],
                             in_data[744],
                             in_data[368],
                             in_data[699],
                             in_data[452]};
    
    wire lut_1364_out = lut_1364_table[lut_1364_select];
    
    generate
    if ( USE_REG ) begin : ff_1364
        reg   lut_1364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1364_ff <= lut_1364_out;
            end
        end
        
        assign out_data[1364] = lut_1364_ff;
    end
    else begin : no_ff_1364
        assign out_data[1364] = lut_1364_out;
    end
    endgenerate
    
    
    
    // LUT : 1365
    wire [63:0] lut_1365_table = 64'b0000000000000000000011110000010100000000000000000000111100001101;
    wire [5:0] lut_1365_select = {
                             in_data[402],
                             in_data[97],
                             in_data[53],
                             in_data[204],
                             in_data[393],
                             in_data[216]};
    
    wire lut_1365_out = lut_1365_table[lut_1365_select];
    
    generate
    if ( USE_REG ) begin : ff_1365
        reg   lut_1365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1365_ff <= lut_1365_out;
            end
        end
        
        assign out_data[1365] = lut_1365_ff;
    end
    else begin : no_ff_1365
        assign out_data[1365] = lut_1365_out;
    end
    endgenerate
    
    
    
    // LUT : 1366
    wire [63:0] lut_1366_table = 64'b1111111011111111111111001111111011111110111111111111110011111000;
    wire [5:0] lut_1366_select = {
                             in_data[728],
                             in_data[496],
                             in_data[118],
                             in_data[509],
                             in_data[371],
                             in_data[747]};
    
    wire lut_1366_out = lut_1366_table[lut_1366_select];
    
    generate
    if ( USE_REG ) begin : ff_1366
        reg   lut_1366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1366_ff <= lut_1366_out;
            end
        end
        
        assign out_data[1366] = lut_1366_ff;
    end
    else begin : no_ff_1366
        assign out_data[1366] = lut_1366_out;
    end
    endgenerate
    
    
    
    // LUT : 1367
    wire [63:0] lut_1367_table = 64'b0000000000000000111111111101111100000000000000001111111011111101;
    wire [5:0] lut_1367_select = {
                             in_data[7],
                             in_data[595],
                             in_data[590],
                             in_data[504],
                             in_data[300],
                             in_data[27]};
    
    wire lut_1367_out = lut_1367_table[lut_1367_select];
    
    generate
    if ( USE_REG ) begin : ff_1367
        reg   lut_1367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1367_ff <= lut_1367_out;
            end
        end
        
        assign out_data[1367] = lut_1367_ff;
    end
    else begin : no_ff_1367
        assign out_data[1367] = lut_1367_out;
    end
    endgenerate
    
    
    
    // LUT : 1368
    wire [63:0] lut_1368_table = 64'b1101111111111111110111111111111101001100010011000100110001001100;
    wire [5:0] lut_1368_select = {
                             in_data[473],
                             in_data[754],
                             in_data[560],
                             in_data[771],
                             in_data[542],
                             in_data[281]};
    
    wire lut_1368_out = lut_1368_table[lut_1368_select];
    
    generate
    if ( USE_REG ) begin : ff_1368
        reg   lut_1368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1368_ff <= lut_1368_out;
            end
        end
        
        assign out_data[1368] = lut_1368_ff;
    end
    else begin : no_ff_1368
        assign out_data[1368] = lut_1368_out;
    end
    endgenerate
    
    
    
    // LUT : 1369
    wire [63:0] lut_1369_table = 64'b0000000000000000000000001111111100000000000000000000000011111111;
    wire [5:0] lut_1369_select = {
                             in_data[670],
                             in_data[369],
                             in_data[330],
                             in_data[2],
                             in_data[697],
                             in_data[325]};
    
    wire lut_1369_out = lut_1369_table[lut_1369_select];
    
    generate
    if ( USE_REG ) begin : ff_1369
        reg   lut_1369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1369_ff <= lut_1369_out;
            end
        end
        
        assign out_data[1369] = lut_1369_ff;
    end
    else begin : no_ff_1369
        assign out_data[1369] = lut_1369_out;
    end
    endgenerate
    
    
    
    // LUT : 1370
    wire [63:0] lut_1370_table = 64'b1111111110111011111111110010001010111011101110111011101100100010;
    wire [5:0] lut_1370_select = {
                             in_data[154],
                             in_data[523],
                             in_data[442],
                             in_data[532],
                             in_data[255],
                             in_data[472]};
    
    wire lut_1370_out = lut_1370_table[lut_1370_select];
    
    generate
    if ( USE_REG ) begin : ff_1370
        reg   lut_1370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1370_ff <= lut_1370_out;
            end
        end
        
        assign out_data[1370] = lut_1370_ff;
    end
    else begin : no_ff_1370
        assign out_data[1370] = lut_1370_out;
    end
    endgenerate
    
    
    
    // LUT : 1371
    wire [63:0] lut_1371_table = 64'b0000000000000000101010101010101000000000000000001010101010101010;
    wire [5:0] lut_1371_select = {
                             in_data[476],
                             in_data[304],
                             in_data[752],
                             in_data[363],
                             in_data[8],
                             in_data[344]};
    
    wire lut_1371_out = lut_1371_table[lut_1371_select];
    
    generate
    if ( USE_REG ) begin : ff_1371
        reg   lut_1371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1371_ff <= lut_1371_out;
            end
        end
        
        assign out_data[1371] = lut_1371_ff;
    end
    else begin : no_ff_1371
        assign out_data[1371] = lut_1371_out;
    end
    endgenerate
    
    
    
    // LUT : 1372
    wire [63:0] lut_1372_table = 64'b0000000000001010000000000000111100000000000010100000000000001011;
    wire [5:0] lut_1372_select = {
                             in_data[478],
                             in_data[475],
                             in_data[581],
                             in_data[153],
                             in_data[6],
                             in_data[412]};
    
    wire lut_1372_out = lut_1372_table[lut_1372_select];
    
    generate
    if ( USE_REG ) begin : ff_1372
        reg   lut_1372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1372_ff <= lut_1372_out;
            end
        end
        
        assign out_data[1372] = lut_1372_ff;
    end
    else begin : no_ff_1372
        assign out_data[1372] = lut_1372_out;
    end
    endgenerate
    
    
    
    // LUT : 1373
    wire [63:0] lut_1373_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1373_select = {
                             in_data[184],
                             in_data[671],
                             in_data[55],
                             in_data[707],
                             in_data[488],
                             in_data[39]};
    
    wire lut_1373_out = lut_1373_table[lut_1373_select];
    
    generate
    if ( USE_REG ) begin : ff_1373
        reg   lut_1373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1373_ff <= lut_1373_out;
            end
        end
        
        assign out_data[1373] = lut_1373_ff;
    end
    else begin : no_ff_1373
        assign out_data[1373] = lut_1373_out;
    end
    endgenerate
    
    
    
    // LUT : 1374
    wire [63:0] lut_1374_table = 64'b0000000000000000000000000000000000000000010101010000000000000100;
    wire [5:0] lut_1374_select = {
                             in_data[593],
                             in_data[319],
                             in_data[770],
                             in_data[591],
                             in_data[701],
                             in_data[635]};
    
    wire lut_1374_out = lut_1374_table[lut_1374_select];
    
    generate
    if ( USE_REG ) begin : ff_1374
        reg   lut_1374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1374_ff <= lut_1374_out;
            end
        end
        
        assign out_data[1374] = lut_1374_ff;
    end
    else begin : no_ff_1374
        assign out_data[1374] = lut_1374_out;
    end
    endgenerate
    
    
    
    // LUT : 1375
    wire [63:0] lut_1375_table = 64'b1111111111101111111111011101010011111111110011001111010111010000;
    wire [5:0] lut_1375_select = {
                             in_data[285],
                             in_data[463],
                             in_data[235],
                             in_data[432],
                             in_data[288],
                             in_data[161]};
    
    wire lut_1375_out = lut_1375_table[lut_1375_select];
    
    generate
    if ( USE_REG ) begin : ff_1375
        reg   lut_1375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1375_ff <= lut_1375_out;
            end
        end
        
        assign out_data[1375] = lut_1375_ff;
    end
    else begin : no_ff_1375
        assign out_data[1375] = lut_1375_out;
    end
    endgenerate
    
    
    
    // LUT : 1376
    wire [63:0] lut_1376_table = 64'b0001001100010011001101110011001100000001000000000001000100000000;
    wire [5:0] lut_1376_select = {
                             in_data[358],
                             in_data[648],
                             in_data[117],
                             in_data[391],
                             in_data[130],
                             in_data[174]};
    
    wire lut_1376_out = lut_1376_table[lut_1376_select];
    
    generate
    if ( USE_REG ) begin : ff_1376
        reg   lut_1376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1376_ff <= lut_1376_out;
            end
        end
        
        assign out_data[1376] = lut_1376_ff;
    end
    else begin : no_ff_1376
        assign out_data[1376] = lut_1376_out;
    end
    endgenerate
    
    
    
    // LUT : 1377
    wire [63:0] lut_1377_table = 64'b0001000000000000000100000000000001110011000000000011001100000000;
    wire [5:0] lut_1377_select = {
                             in_data[668],
                             in_data[30],
                             in_data[370],
                             in_data[779],
                             in_data[445],
                             in_data[88]};
    
    wire lut_1377_out = lut_1377_table[lut_1377_select];
    
    generate
    if ( USE_REG ) begin : ff_1377
        reg   lut_1377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1377_ff <= lut_1377_out;
            end
        end
        
        assign out_data[1377] = lut_1377_ff;
    end
    else begin : no_ff_1377
        assign out_data[1377] = lut_1377_out;
    end
    endgenerate
    
    
    
    // LUT : 1378
    wire [63:0] lut_1378_table = 64'b1111001111110011110100001101000111110111111101111101000011010001;
    wire [5:0] lut_1378_select = {
                             in_data[317],
                             in_data[481],
                             in_data[748],
                             in_data[547],
                             in_data[230],
                             in_data[406]};
    
    wire lut_1378_out = lut_1378_table[lut_1378_select];
    
    generate
    if ( USE_REG ) begin : ff_1378
        reg   lut_1378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1378_ff <= lut_1378_out;
            end
        end
        
        assign out_data[1378] = lut_1378_ff;
    end
    else begin : no_ff_1378
        assign out_data[1378] = lut_1378_out;
    end
    endgenerate
    
    
    
    // LUT : 1379
    wire [63:0] lut_1379_table = 64'b1010111111111111101011111101111110101111000001011010111100000101;
    wire [5:0] lut_1379_select = {
                             in_data[233],
                             in_data[727],
                             in_data[208],
                             in_data[221],
                             in_data[725],
                             in_data[297]};
    
    wire lut_1379_out = lut_1379_table[lut_1379_select];
    
    generate
    if ( USE_REG ) begin : ff_1379
        reg   lut_1379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1379_ff <= lut_1379_out;
            end
        end
        
        assign out_data[1379] = lut_1379_ff;
    end
    else begin : no_ff_1379
        assign out_data[1379] = lut_1379_out;
    end
    endgenerate
    
    
    
    // LUT : 1380
    wire [63:0] lut_1380_table = 64'b0011110010111100101111001011110011111100111111001011110010111100;
    wire [5:0] lut_1380_select = {
                             in_data[195],
                             in_data[759],
                             in_data[503],
                             in_data[551],
                             in_data[213],
                             in_data[41]};
    
    wire lut_1380_out = lut_1380_table[lut_1380_select];
    
    generate
    if ( USE_REG ) begin : ff_1380
        reg   lut_1380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1380_ff <= lut_1380_out;
            end
        end
        
        assign out_data[1380] = lut_1380_ff;
    end
    else begin : no_ff_1380
        assign out_data[1380] = lut_1380_out;
    end
    endgenerate
    
    
    
    // LUT : 1381
    wire [63:0] lut_1381_table = 64'b1111111111111111111111110000000011111111111111111111111100000000;
    wire [5:0] lut_1381_select = {
                             in_data[757],
                             in_data[400],
                             in_data[693],
                             in_data[470],
                             in_data[43],
                             in_data[225]};
    
    wire lut_1381_out = lut_1381_table[lut_1381_select];
    
    generate
    if ( USE_REG ) begin : ff_1381
        reg   lut_1381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1381_ff <= lut_1381_out;
            end
        end
        
        assign out_data[1381] = lut_1381_ff;
    end
    else begin : no_ff_1381
        assign out_data[1381] = lut_1381_out;
    end
    endgenerate
    
    
    
    // LUT : 1382
    wire [63:0] lut_1382_table = 64'b0000100010001000000000000000000000000000100011001100110010111011;
    wire [5:0] lut_1382_select = {
                             in_data[157],
                             in_data[623],
                             in_data[539],
                             in_data[756],
                             in_data[155],
                             in_data[681]};
    
    wire lut_1382_out = lut_1382_table[lut_1382_select];
    
    generate
    if ( USE_REG ) begin : ff_1382
        reg   lut_1382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1382_ff <= lut_1382_out;
            end
        end
        
        assign out_data[1382] = lut_1382_ff;
    end
    else begin : no_ff_1382
        assign out_data[1382] = lut_1382_out;
    end
    endgenerate
    
    
    
    // LUT : 1383
    wire [63:0] lut_1383_table = 64'b0000000000001111000011100000111100001000000011110000111000001111;
    wire [5:0] lut_1383_select = {
                             in_data[589],
                             in_data[489],
                             in_data[490],
                             in_data[535],
                             in_data[376],
                             in_data[666]};
    
    wire lut_1383_out = lut_1383_table[lut_1383_select];
    
    generate
    if ( USE_REG ) begin : ff_1383
        reg   lut_1383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1383_ff <= lut_1383_out;
            end
        end
        
        assign out_data[1383] = lut_1383_ff;
    end
    else begin : no_ff_1383
        assign out_data[1383] = lut_1383_out;
    end
    endgenerate
    
    
    
    // LUT : 1384
    wire [63:0] lut_1384_table = 64'b0000000000111111000000000011111100000000001111110000000000111111;
    wire [5:0] lut_1384_select = {
                             in_data[421],
                             in_data[38],
                             in_data[525],
                             in_data[544],
                             in_data[415],
                             in_data[114]};
    
    wire lut_1384_out = lut_1384_table[lut_1384_select];
    
    generate
    if ( USE_REG ) begin : ff_1384
        reg   lut_1384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1384_ff <= lut_1384_out;
            end
        end
        
        assign out_data[1384] = lut_1384_ff;
    end
    else begin : no_ff_1384
        assign out_data[1384] = lut_1384_out;
    end
    endgenerate
    
    
    
    // LUT : 1385
    wire [63:0] lut_1385_table = 64'b0000000000000000000011110010111100000000000000000000111100011111;
    wire [5:0] lut_1385_select = {
                             in_data[494],
                             in_data[456],
                             in_data[610],
                             in_data[411],
                             in_data[690],
                             in_data[163]};
    
    wire lut_1385_out = lut_1385_table[lut_1385_select];
    
    generate
    if ( USE_REG ) begin : ff_1385
        reg   lut_1385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1385_ff <= lut_1385_out;
            end
        end
        
        assign out_data[1385] = lut_1385_ff;
    end
    else begin : no_ff_1385
        assign out_data[1385] = lut_1385_out;
    end
    endgenerate
    
    
    
    // LUT : 1386
    wire [63:0] lut_1386_table = 64'b1011101110111011101110111011101110111011101110111011101110111011;
    wire [5:0] lut_1386_select = {
                             in_data[26],
                             in_data[110],
                             in_data[528],
                             in_data[588],
                             in_data[429],
                             in_data[74]};
    
    wire lut_1386_out = lut_1386_table[lut_1386_select];
    
    generate
    if ( USE_REG ) begin : ff_1386
        reg   lut_1386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1386_ff <= lut_1386_out;
            end
        end
        
        assign out_data[1386] = lut_1386_ff;
    end
    else begin : no_ff_1386
        assign out_data[1386] = lut_1386_out;
    end
    endgenerate
    
    
    
    // LUT : 1387
    wire [63:0] lut_1387_table = 64'b1100110011001100110011001100110011111111111111111111111111111111;
    wire [5:0] lut_1387_select = {
                             in_data[243],
                             in_data[64],
                             in_data[52],
                             in_data[5],
                             in_data[202],
                             in_data[559]};
    
    wire lut_1387_out = lut_1387_table[lut_1387_select];
    
    generate
    if ( USE_REG ) begin : ff_1387
        reg   lut_1387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1387_ff <= lut_1387_out;
            end
        end
        
        assign out_data[1387] = lut_1387_ff;
    end
    else begin : no_ff_1387
        assign out_data[1387] = lut_1387_out;
    end
    endgenerate
    
    
    
    // LUT : 1388
    wire [63:0] lut_1388_table = 64'b0000000000000000000000000000000011111111111011111111111111001111;
    wire [5:0] lut_1388_select = {
                             in_data[180],
                             in_data[256],
                             in_data[107],
                             in_data[278],
                             in_data[314],
                             in_data[694]};
    
    wire lut_1388_out = lut_1388_table[lut_1388_select];
    
    generate
    if ( USE_REG ) begin : ff_1388
        reg   lut_1388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1388_ff <= lut_1388_out;
            end
        end
        
        assign out_data[1388] = lut_1388_ff;
    end
    else begin : no_ff_1388
        assign out_data[1388] = lut_1388_out;
    end
    endgenerate
    
    
    
    // LUT : 1389
    wire [63:0] lut_1389_table = 64'b0000000000000000000001010000010100000000000000000000111100001111;
    wire [5:0] lut_1389_select = {
                             in_data[331],
                             in_data[373],
                             in_data[166],
                             in_data[580],
                             in_data[251],
                             in_data[482]};
    
    wire lut_1389_out = lut_1389_table[lut_1389_select];
    
    generate
    if ( USE_REG ) begin : ff_1389
        reg   lut_1389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1389_ff <= lut_1389_out;
            end
        end
        
        assign out_data[1389] = lut_1389_ff;
    end
    else begin : no_ff_1389
        assign out_data[1389] = lut_1389_out;
    end
    endgenerate
    
    
    
    // LUT : 1390
    wire [63:0] lut_1390_table = 64'b1111111111111111000011100000111111111111111111110000111100001111;
    wire [5:0] lut_1390_select = {
                             in_data[58],
                             in_data[289],
                             in_data[731],
                             in_data[522],
                             in_data[274],
                             in_data[215]};
    
    wire lut_1390_out = lut_1390_table[lut_1390_select];
    
    generate
    if ( USE_REG ) begin : ff_1390
        reg   lut_1390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1390_ff <= lut_1390_out;
            end
        end
        
        assign out_data[1390] = lut_1390_ff;
    end
    else begin : no_ff_1390
        assign out_data[1390] = lut_1390_out;
    end
    endgenerate
    
    
    
    // LUT : 1391
    wire [63:0] lut_1391_table = 64'b0011011100110111001101110011001100110011000100110001000100010011;
    wire [5:0] lut_1391_select = {
                             in_data[571],
                             in_data[87],
                             in_data[422],
                             in_data[737],
                             in_data[438],
                             in_data[647]};
    
    wire lut_1391_out = lut_1391_table[lut_1391_select];
    
    generate
    if ( USE_REG ) begin : ff_1391
        reg   lut_1391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1391_ff <= lut_1391_out;
            end
        end
        
        assign out_data[1391] = lut_1391_ff;
    end
    else begin : no_ff_1391
        assign out_data[1391] = lut_1391_out;
    end
    endgenerate
    
    
    
    // LUT : 1392
    wire [63:0] lut_1392_table = 64'b0000000000000000000000000000000000000000000000001111111111111111;
    wire [5:0] lut_1392_select = {
                             in_data[321],
                             in_data[390],
                             in_data[776],
                             in_data[751],
                             in_data[112],
                             in_data[15]};
    
    wire lut_1392_out = lut_1392_table[lut_1392_select];
    
    generate
    if ( USE_REG ) begin : ff_1392
        reg   lut_1392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1392_ff <= lut_1392_out;
            end
        end
        
        assign out_data[1392] = lut_1392_ff;
    end
    else begin : no_ff_1392
        assign out_data[1392] = lut_1392_out;
    end
    endgenerate
    
    
    
    // LUT : 1393
    wire [63:0] lut_1393_table = 64'b1111111111110000111100000000000011110000111100001111000011110000;
    wire [5:0] lut_1393_select = {
                             in_data[431],
                             in_data[657],
                             in_data[257],
                             in_data[439],
                             in_data[782],
                             in_data[614]};
    
    wire lut_1393_out = lut_1393_table[lut_1393_select];
    
    generate
    if ( USE_REG ) begin : ff_1393
        reg   lut_1393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1393_ff <= lut_1393_out;
            end
        end
        
        assign out_data[1393] = lut_1393_ff;
    end
    else begin : no_ff_1393
        assign out_data[1393] = lut_1393_out;
    end
    endgenerate
    
    
    
    // LUT : 1394
    wire [63:0] lut_1394_table = 64'b1100110011001100100011001100110011001100110011000000110011001100;
    wire [5:0] lut_1394_select = {
                             in_data[394],
                             in_data[70],
                             in_data[695],
                             in_data[565],
                             in_data[469],
                             in_data[333]};
    
    wire lut_1394_out = lut_1394_table[lut_1394_select];
    
    generate
    if ( USE_REG ) begin : ff_1394
        reg   lut_1394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1394_ff <= lut_1394_out;
            end
        end
        
        assign out_data[1394] = lut_1394_ff;
    end
    else begin : no_ff_1394
        assign out_data[1394] = lut_1394_out;
    end
    endgenerate
    
    
    
    // LUT : 1395
    wire [63:0] lut_1395_table = 64'b1011101111111111111111111111111100000010101110111100110001010101;
    wire [5:0] lut_1395_select = {
                             in_data[340],
                             in_data[577],
                             in_data[385],
                             in_data[618],
                             in_data[655],
                             in_data[234]};
    
    wire lut_1395_out = lut_1395_table[lut_1395_select];
    
    generate
    if ( USE_REG ) begin : ff_1395
        reg   lut_1395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1395_ff <= lut_1395_out;
            end
        end
        
        assign out_data[1395] = lut_1395_ff;
    end
    else begin : no_ff_1395
        assign out_data[1395] = lut_1395_out;
    end
    endgenerate
    
    
    
    // LUT : 1396
    wire [63:0] lut_1396_table = 64'b0001000000000000111100001111000111110000010100001111000111111101;
    wire [5:0] lut_1396_select = {
                             in_data[461],
                             in_data[650],
                             in_data[594],
                             in_data[247],
                             in_data[596],
                             in_data[497]};
    
    wire lut_1396_out = lut_1396_table[lut_1396_select];
    
    generate
    if ( USE_REG ) begin : ff_1396
        reg   lut_1396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1396_ff <= lut_1396_out;
            end
        end
        
        assign out_data[1396] = lut_1396_ff;
    end
    else begin : no_ff_1396
        assign out_data[1396] = lut_1396_out;
    end
    endgenerate
    
    
    
    // LUT : 1397
    wire [63:0] lut_1397_table = 64'b0000010100000101000001010000010100000101000001010000010100000101;
    wire [5:0] lut_1397_select = {
                             in_data[569],
                             in_data[45],
                             in_data[505],
                             in_data[453],
                             in_data[334],
                             in_data[454]};
    
    wire lut_1397_out = lut_1397_table[lut_1397_select];
    
    generate
    if ( USE_REG ) begin : ff_1397
        reg   lut_1397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1397_ff <= lut_1397_out;
            end
        end
        
        assign out_data[1397] = lut_1397_ff;
    end
    else begin : no_ff_1397
        assign out_data[1397] = lut_1397_out;
    end
    endgenerate
    
    
    
    // LUT : 1398
    wire [63:0] lut_1398_table = 64'b1100110111001101110011011100110011001101010001001100110100000100;
    wire [5:0] lut_1398_select = {
                             in_data[769],
                             in_data[774],
                             in_data[708],
                             in_data[276],
                             in_data[495],
                             in_data[567]};
    
    wire lut_1398_out = lut_1398_table[lut_1398_select];
    
    generate
    if ( USE_REG ) begin : ff_1398
        reg   lut_1398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1398_ff <= lut_1398_out;
            end
        end
        
        assign out_data[1398] = lut_1398_ff;
    end
    else begin : no_ff_1398
        assign out_data[1398] = lut_1398_out;
    end
    endgenerate
    
    
    
    // LUT : 1399
    wire [63:0] lut_1399_table = 64'b1111111111001100110011000000000011111111111111111111111111111100;
    wire [5:0] lut_1399_select = {
                             in_data[483],
                             in_data[518],
                             in_data[203],
                             in_data[682],
                             in_data[246],
                             in_data[132]};
    
    wire lut_1399_out = lut_1399_table[lut_1399_select];
    
    generate
    if ( USE_REG ) begin : ff_1399
        reg   lut_1399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1399_ff <= lut_1399_out;
            end
        end
        
        assign out_data[1399] = lut_1399_ff;
    end
    else begin : no_ff_1399
        assign out_data[1399] = lut_1399_out;
    end
    endgenerate
    
    
    
    // LUT : 1400
    wire [63:0] lut_1400_table = 64'b0000000011001100000000001100110000000000111111111100000011111111;
    wire [5:0] lut_1400_select = {
                             in_data[378],
                             in_data[691],
                             in_data[137],
                             in_data[738],
                             in_data[67],
                             in_data[778]};
    
    wire lut_1400_out = lut_1400_table[lut_1400_select];
    
    generate
    if ( USE_REG ) begin : ff_1400
        reg   lut_1400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1400_ff <= lut_1400_out;
            end
        end
        
        assign out_data[1400] = lut_1400_ff;
    end
    else begin : no_ff_1400
        assign out_data[1400] = lut_1400_out;
    end
    endgenerate
    
    
    
    // LUT : 1401
    wire [63:0] lut_1401_table = 64'b1111111111111111111111111111111111101100101010000100010010001110;
    wire [5:0] lut_1401_select = {
                             in_data[295],
                             in_data[409],
                             in_data[713],
                             in_data[741],
                             in_data[677],
                             in_data[654]};
    
    wire lut_1401_out = lut_1401_table[lut_1401_select];
    
    generate
    if ( USE_REG ) begin : ff_1401
        reg   lut_1401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1401_ff <= lut_1401_out;
            end
        end
        
        assign out_data[1401] = lut_1401_ff;
    end
    else begin : no_ff_1401
        assign out_data[1401] = lut_1401_out;
    end
    endgenerate
    
    
    
    // LUT : 1402
    wire [63:0] lut_1402_table = 64'b0000000000000000001111110011111100000000000000000000111100001111;
    wire [5:0] lut_1402_select = {
                             in_data[236],
                             in_data[659],
                             in_data[730],
                             in_data[266],
                             in_data[265],
                             in_data[11]};
    
    wire lut_1402_out = lut_1402_table[lut_1402_select];
    
    generate
    if ( USE_REG ) begin : ff_1402
        reg   lut_1402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1402_ff <= lut_1402_out;
            end
        end
        
        assign out_data[1402] = lut_1402_ff;
    end
    else begin : no_ff_1402
        assign out_data[1402] = lut_1402_out;
    end
    endgenerate
    
    
    
    // LUT : 1403
    wire [63:0] lut_1403_table = 64'b0000000000000000000000000000111100000000001011110000000011111111;
    wire [5:0] lut_1403_select = {
                             in_data[121],
                             in_data[709],
                             in_data[575],
                             in_data[149],
                             in_data[566],
                             in_data[606]};
    
    wire lut_1403_out = lut_1403_table[lut_1403_select];
    
    generate
    if ( USE_REG ) begin : ff_1403
        reg   lut_1403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1403_ff <= lut_1403_out;
            end
        end
        
        assign out_data[1403] = lut_1403_ff;
    end
    else begin : no_ff_1403
        assign out_data[1403] = lut_1403_out;
    end
    endgenerate
    
    
    
    // LUT : 1404
    wire [63:0] lut_1404_table = 64'b0010000000100000111100111011001100110011001100111011001100110011;
    wire [5:0] lut_1404_select = {
                             in_data[239],
                             in_data[187],
                             in_data[227],
                             in_data[468],
                             in_data[181],
                             in_data[228]};
    
    wire lut_1404_out = lut_1404_table[lut_1404_select];
    
    generate
    if ( USE_REG ) begin : ff_1404
        reg   lut_1404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1404_ff <= lut_1404_out;
            end
        end
        
        assign out_data[1404] = lut_1404_ff;
    end
    else begin : no_ff_1404
        assign out_data[1404] = lut_1404_out;
    end
    endgenerate
    
    
    
    // LUT : 1405
    wire [63:0] lut_1405_table = 64'b0000000000000010000000000000001000000000000000010000000000000001;
    wire [5:0] lut_1405_select = {
                             in_data[617],
                             in_data[140],
                             in_data[102],
                             in_data[108],
                             in_data[703],
                             in_data[755]};
    
    wire lut_1405_out = lut_1405_table[lut_1405_select];
    
    generate
    if ( USE_REG ) begin : ff_1405
        reg   lut_1405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1405_ff <= lut_1405_out;
            end
        end
        
        assign out_data[1405] = lut_1405_ff;
    end
    else begin : no_ff_1405
        assign out_data[1405] = lut_1405_out;
    end
    endgenerate
    
    
    
    // LUT : 1406
    wire [63:0] lut_1406_table = 64'b1100110011101100110011001110110011111100111111101111110011111111;
    wire [5:0] lut_1406_select = {
                             in_data[527],
                             in_data[767],
                             in_data[179],
                             in_data[162],
                             in_data[679],
                             in_data[717]};
    
    wire lut_1406_out = lut_1406_table[lut_1406_select];
    
    generate
    if ( USE_REG ) begin : ff_1406
        reg   lut_1406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1406_ff <= lut_1406_out;
            end
        end
        
        assign out_data[1406] = lut_1406_ff;
    end
    else begin : no_ff_1406
        assign out_data[1406] = lut_1406_out;
    end
    endgenerate
    
    
    
    // LUT : 1407
    wire [63:0] lut_1407_table = 64'b0000000000000000010100000101000000000000000000000101000001010001;
    wire [5:0] lut_1407_select = {
                             in_data[361],
                             in_data[578],
                             in_data[530],
                             in_data[346],
                             in_data[457],
                             in_data[636]};
    
    wire lut_1407_out = lut_1407_table[lut_1407_select];
    
    generate
    if ( USE_REG ) begin : ff_1407
        reg   lut_1407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1407_ff <= lut_1407_out;
            end
        end
        
        assign out_data[1407] = lut_1407_ff;
    end
    else begin : no_ff_1407
        assign out_data[1407] = lut_1407_out;
    end
    endgenerate
    
    
    
    // LUT : 1408
    wire [63:0] lut_1408_table = 64'b0000000000000000000000000000000000000001000101010000000001000101;
    wire [5:0] lut_1408_select = {
                             in_data[582],
                             in_data[602],
                             in_data[190],
                             in_data[619],
                             in_data[122],
                             in_data[404]};
    
    wire lut_1408_out = lut_1408_table[lut_1408_select];
    
    generate
    if ( USE_REG ) begin : ff_1408
        reg   lut_1408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1408_ff <= lut_1408_out;
            end
        end
        
        assign out_data[1408] = lut_1408_ff;
    end
    else begin : no_ff_1408
        assign out_data[1408] = lut_1408_out;
    end
    endgenerate
    
    
    
    // LUT : 1409
    wire [63:0] lut_1409_table = 64'b1111111111111111000011100000000011111111111111110000111000000000;
    wire [5:0] lut_1409_select = {
                             in_data[702],
                             in_data[377],
                             in_data[76],
                             in_data[170],
                             in_data[51],
                             in_data[533]};
    
    wire lut_1409_out = lut_1409_table[lut_1409_select];
    
    generate
    if ( USE_REG ) begin : ff_1409
        reg   lut_1409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1409_ff <= lut_1409_out;
            end
        end
        
        assign out_data[1409] = lut_1409_ff;
    end
    else begin : no_ff_1409
        assign out_data[1409] = lut_1409_out;
    end
    endgenerate
    
    
    
    // LUT : 1410
    wire [63:0] lut_1410_table = 64'b0000000011111111000000000000111100000000111111110000000000001111;
    wire [5:0] lut_1410_select = {
                             in_data[169],
                             in_data[396],
                             in_data[430],
                             in_data[397],
                             in_data[447],
                             in_data[57]};
    
    wire lut_1410_out = lut_1410_table[lut_1410_select];
    
    generate
    if ( USE_REG ) begin : ff_1410
        reg   lut_1410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1410_ff <= lut_1410_out;
            end
        end
        
        assign out_data[1410] = lut_1410_ff;
    end
    else begin : no_ff_1410
        assign out_data[1410] = lut_1410_out;
    end
    endgenerate
    
    
    
    // LUT : 1411
    wire [63:0] lut_1411_table = 64'b1111111111111111111111111111111100000000001111110000000000000000;
    wire [5:0] lut_1411_select = {
                             in_data[275],
                             in_data[405],
                             in_data[408],
                             in_data[364],
                             in_data[135],
                             in_data[24]};
    
    wire lut_1411_out = lut_1411_table[lut_1411_select];
    
    generate
    if ( USE_REG ) begin : ff_1411
        reg   lut_1411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1411_ff <= lut_1411_out;
            end
        end
        
        assign out_data[1411] = lut_1411_ff;
    end
    else begin : no_ff_1411
        assign out_data[1411] = lut_1411_out;
    end
    endgenerate
    
    
    
    // LUT : 1412
    wire [63:0] lut_1412_table = 64'b1010101111111111111111111111111110001000100010001011101110001010;
    wire [5:0] lut_1412_select = {
                             in_data[220],
                             in_data[462],
                             in_data[632],
                             in_data[446],
                             in_data[286],
                             in_data[426]};
    
    wire lut_1412_out = lut_1412_table[lut_1412_select];
    
    generate
    if ( USE_REG ) begin : ff_1412
        reg   lut_1412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1412_ff <= lut_1412_out;
            end
        end
        
        assign out_data[1412] = lut_1412_ff;
    end
    else begin : no_ff_1412
        assign out_data[1412] = lut_1412_out;
    end
    endgenerate
    
    
    
    // LUT : 1413
    wire [63:0] lut_1413_table = 64'b0000010100000101000001010000010100000000000000000000000000000000;
    wire [5:0] lut_1413_select = {
                             in_data[441],
                             in_data[60],
                             in_data[34],
                             in_data[315],
                             in_data[14],
                             in_data[665]};
    
    wire lut_1413_out = lut_1413_table[lut_1413_select];
    
    generate
    if ( USE_REG ) begin : ff_1413
        reg   lut_1413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1413_ff <= lut_1413_out;
            end
        end
        
        assign out_data[1413] = lut_1413_ff;
    end
    else begin : no_ff_1413
        assign out_data[1413] = lut_1413_out;
    end
    endgenerate
    
    
    
    // LUT : 1414
    wire [63:0] lut_1414_table = 64'b0000000100000000111111111111111100010000000100001111010111110101;
    wire [5:0] lut_1414_select = {
                             in_data[205],
                             in_data[382],
                             in_data[66],
                             in_data[126],
                             in_data[29],
                             in_data[328]};
    
    wire lut_1414_out = lut_1414_table[lut_1414_select];
    
    generate
    if ( USE_REG ) begin : ff_1414
        reg   lut_1414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1414_ff <= lut_1414_out;
            end
        end
        
        assign out_data[1414] = lut_1414_ff;
    end
    else begin : no_ff_1414
        assign out_data[1414] = lut_1414_out;
    end
    endgenerate
    
    
    
    // LUT : 1415
    wire [63:0] lut_1415_table = 64'b1111111111111111000000110000000011111111111111110000001100000000;
    wire [5:0] lut_1415_select = {
                             in_data[23],
                             in_data[326],
                             in_data[277],
                             in_data[658],
                             in_data[188],
                             in_data[477]};
    
    wire lut_1415_out = lut_1415_table[lut_1415_select];
    
    generate
    if ( USE_REG ) begin : ff_1415
        reg   lut_1415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1415_ff <= lut_1415_out;
            end
        end
        
        assign out_data[1415] = lut_1415_ff;
    end
    else begin : no_ff_1415
        assign out_data[1415] = lut_1415_out;
    end
    endgenerate
    
    
    
    // LUT : 1416
    wire [63:0] lut_1416_table = 64'b0000000000000000010101010101010100000100000001000101010101010101;
    wire [5:0] lut_1416_select = {
                             in_data[419],
                             in_data[241],
                             in_data[534],
                             in_data[271],
                             in_data[10],
                             in_data[711]};
    
    wire lut_1416_out = lut_1416_table[lut_1416_select];
    
    generate
    if ( USE_REG ) begin : ff_1416
        reg   lut_1416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1416_ff <= lut_1416_out;
            end
        end
        
        assign out_data[1416] = lut_1416_ff;
    end
    else begin : no_ff_1416
        assign out_data[1416] = lut_1416_out;
    end
    endgenerate
    
    
    
    // LUT : 1417
    wire [63:0] lut_1417_table = 64'b0000000000000000000000000000000010111011101110111010101110101011;
    wire [5:0] lut_1417_select = {
                             in_data[159],
                             in_data[353],
                             in_data[698],
                             in_data[44],
                             in_data[718],
                             in_data[395]};
    
    wire lut_1417_out = lut_1417_table[lut_1417_select];
    
    generate
    if ( USE_REG ) begin : ff_1417
        reg   lut_1417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1417_ff <= lut_1417_out;
            end
        end
        
        assign out_data[1417] = lut_1417_ff;
    end
    else begin : no_ff_1417
        assign out_data[1417] = lut_1417_out;
    end
    endgenerate
    
    
    
    // LUT : 1418
    wire [63:0] lut_1418_table = 64'b0000000000000000000000000000000011011111010111111101111101011111;
    wire [5:0] lut_1418_select = {
                             in_data[656],
                             in_data[674],
                             in_data[519],
                             in_data[232],
                             in_data[337],
                             in_data[296]};
    
    wire lut_1418_out = lut_1418_table[lut_1418_select];
    
    generate
    if ( USE_REG ) begin : ff_1418
        reg   lut_1418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1418_ff <= lut_1418_out;
            end
        end
        
        assign out_data[1418] = lut_1418_ff;
    end
    else begin : no_ff_1418
        assign out_data[1418] = lut_1418_out;
    end
    endgenerate
    
    
    
    // LUT : 1419
    wire [63:0] lut_1419_table = 64'b1111111111111100111111101111111011111111111111111111110011111100;
    wire [5:0] lut_1419_select = {
                             in_data[631],
                             in_data[499],
                             in_data[620],
                             in_data[305],
                             in_data[434],
                             in_data[634]};
    
    wire lut_1419_out = lut_1419_table[lut_1419_select];
    
    generate
    if ( USE_REG ) begin : ff_1419
        reg   lut_1419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1419_ff <= lut_1419_out;
            end
        end
        
        assign out_data[1419] = lut_1419_ff;
    end
    else begin : no_ff_1419
        assign out_data[1419] = lut_1419_out;
    end
    endgenerate
    
    
    
    // LUT : 1420
    wire [63:0] lut_1420_table = 64'b0000000000000000010101010101010100000000000000000101010101010101;
    wire [5:0] lut_1420_select = {
                             in_data[733],
                             in_data[359],
                             in_data[766],
                             in_data[63],
                             in_data[3],
                             in_data[301]};
    
    wire lut_1420_out = lut_1420_table[lut_1420_select];
    
    generate
    if ( USE_REG ) begin : ff_1420
        reg   lut_1420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1420_ff <= lut_1420_out;
            end
        end
        
        assign out_data[1420] = lut_1420_ff;
    end
    else begin : no_ff_1420
        assign out_data[1420] = lut_1420_out;
    end
    endgenerate
    
    
    
    // LUT : 1421
    wire [63:0] lut_1421_table = 64'b0000000000111111000000000011111100000000001111110000000000000011;
    wire [5:0] lut_1421_select = {
                             in_data[194],
                             in_data[258],
                             in_data[651],
                             in_data[283],
                             in_data[436],
                             in_data[17]};
    
    wire lut_1421_out = lut_1421_table[lut_1421_select];
    
    generate
    if ( USE_REG ) begin : ff_1421
        reg   lut_1421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1421_ff <= lut_1421_out;
            end
        end
        
        assign out_data[1421] = lut_1421_ff;
    end
    else begin : no_ff_1421
        assign out_data[1421] = lut_1421_out;
    end
    endgenerate
    
    
    
    // LUT : 1422
    wire [63:0] lut_1422_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1422_select = {
                             in_data[327],
                             in_data[585],
                             in_data[253],
                             in_data[360],
                             in_data[604],
                             in_data[22]};
    
    wire lut_1422_out = lut_1422_table[lut_1422_select];
    
    generate
    if ( USE_REG ) begin : ff_1422
        reg   lut_1422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1422_ff <= lut_1422_out;
            end
        end
        
        assign out_data[1422] = lut_1422_ff;
    end
    else begin : no_ff_1422
        assign out_data[1422] = lut_1422_out;
    end
    endgenerate
    
    
    
    // LUT : 1423
    wire [63:0] lut_1423_table = 64'b0100110001000100110011001100110011001100110011001111111111001100;
    wire [5:0] lut_1423_select = {
                             in_data[345],
                             in_data[423],
                             in_data[240],
                             in_data[696],
                             in_data[264],
                             in_data[724]};
    
    wire lut_1423_out = lut_1423_table[lut_1423_select];
    
    generate
    if ( USE_REG ) begin : ff_1423
        reg   lut_1423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1423_ff <= lut_1423_out;
            end
        end
        
        assign out_data[1423] = lut_1423_ff;
    end
    else begin : no_ff_1423
        assign out_data[1423] = lut_1423_out;
    end
    endgenerate
    
    
    
    // LUT : 1424
    wire [63:0] lut_1424_table = 64'b0100010000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1424_select = {
                             in_data[550],
                             in_data[764],
                             in_data[1],
                             in_data[12],
                             in_data[47],
                             in_data[603]};
    
    wire lut_1424_out = lut_1424_table[lut_1424_select];
    
    generate
    if ( USE_REG ) begin : ff_1424
        reg   lut_1424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1424_ff <= lut_1424_out;
            end
        end
        
        assign out_data[1424] = lut_1424_ff;
    end
    else begin : no_ff_1424
        assign out_data[1424] = lut_1424_out;
    end
    endgenerate
    
    
    
    // LUT : 1425
    wire [63:0] lut_1425_table = 64'b1111111111111111111111111111111100100000101000001010101010101010;
    wire [5:0] lut_1425_select = {
                             in_data[298],
                             in_data[127],
                             in_data[336],
                             in_data[366],
                             in_data[750],
                             in_data[417]};
    
    wire lut_1425_out = lut_1425_table[lut_1425_select];
    
    generate
    if ( USE_REG ) begin : ff_1425
        reg   lut_1425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1425_ff <= lut_1425_out;
            end
        end
        
        assign out_data[1425] = lut_1425_ff;
    end
    else begin : no_ff_1425
        assign out_data[1425] = lut_1425_out;
    end
    endgenerate
    
    
    
    // LUT : 1426
    wire [63:0] lut_1426_table = 64'b0000000001000100010101010101010101010101010101010101010101010101;
    wire [5:0] lut_1426_select = {
                             in_data[173],
                             in_data[428],
                             in_data[451],
                             in_data[311],
                             in_data[418],
                             in_data[435]};
    
    wire lut_1426_out = lut_1426_table[lut_1426_select];
    
    generate
    if ( USE_REG ) begin : ff_1426
        reg   lut_1426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1426_ff <= lut_1426_out;
            end
        end
        
        assign out_data[1426] = lut_1426_ff;
    end
    else begin : no_ff_1426
        assign out_data[1426] = lut_1426_out;
    end
    endgenerate
    
    
    
    // LUT : 1427
    wire [63:0] lut_1427_table = 64'b0000110000001100000001000000110000001100000011000000110000001100;
    wire [5:0] lut_1427_select = {
                             in_data[21],
                             in_data[62],
                             in_data[104],
                             in_data[248],
                             in_data[270],
                             in_data[524]};
    
    wire lut_1427_out = lut_1427_table[lut_1427_select];
    
    generate
    if ( USE_REG ) begin : ff_1427
        reg   lut_1427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1427_ff <= lut_1427_out;
            end
        end
        
        assign out_data[1427] = lut_1427_ff;
    end
    else begin : no_ff_1427
        assign out_data[1427] = lut_1427_out;
    end
    endgenerate
    
    
    
    // LUT : 1428
    wire [63:0] lut_1428_table = 64'b1101101011011010111110111111101000010001000100000101000100010001;
    wire [5:0] lut_1428_select = {
                             in_data[440],
                             in_data[742],
                             in_data[736],
                             in_data[347],
                             in_data[350],
                             in_data[433]};
    
    wire lut_1428_out = lut_1428_table[lut_1428_select];
    
    generate
    if ( USE_REG ) begin : ff_1428
        reg   lut_1428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1428_ff <= lut_1428_out;
            end
        end
        
        assign out_data[1428] = lut_1428_ff;
    end
    else begin : no_ff_1428
        assign out_data[1428] = lut_1428_out;
    end
    endgenerate
    
    
    
    // LUT : 1429
    wire [63:0] lut_1429_table = 64'b0111111111111111000000000000000000000000010001000000000001000100;
    wire [5:0] lut_1429_select = {
                             in_data[546],
                             in_data[491],
                             in_data[316],
                             in_data[502],
                             in_data[545],
                             in_data[201]};
    
    wire lut_1429_out = lut_1429_table[lut_1429_select];
    
    generate
    if ( USE_REG ) begin : ff_1429
        reg   lut_1429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1429_ff <= lut_1429_out;
            end
        end
        
        assign out_data[1429] = lut_1429_ff;
    end
    else begin : no_ff_1429
        assign out_data[1429] = lut_1429_out;
    end
    endgenerate
    
    
    
    // LUT : 1430
    wire [63:0] lut_1430_table = 64'b1111111111111111111111111111111100000000000000000011000100110000;
    wire [5:0] lut_1430_select = {
                             in_data[245],
                             in_data[399],
                             in_data[31],
                             in_data[749],
                             in_data[493],
                             in_data[91]};
    
    wire lut_1430_out = lut_1430_table[lut_1430_select];
    
    generate
    if ( USE_REG ) begin : ff_1430
        reg   lut_1430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1430_ff <= lut_1430_out;
            end
        end
        
        assign out_data[1430] = lut_1430_ff;
    end
    else begin : no_ff_1430
        assign out_data[1430] = lut_1430_out;
    end
    endgenerate
    
    
    
    // LUT : 1431
    wire [63:0] lut_1431_table = 64'b1100111100001111110011110000111100000100000011110000010000001111;
    wire [5:0] lut_1431_select = {
                             in_data[654],
                             in_data[755],
                             in_data[522],
                             in_data[487],
                             in_data[736],
                             in_data[204]};
    
    wire lut_1431_out = lut_1431_table[lut_1431_select];
    
    generate
    if ( USE_REG ) begin : ff_1431
        reg   lut_1431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1431_ff <= lut_1431_out;
            end
        end
        
        assign out_data[1431] = lut_1431_ff;
    end
    else begin : no_ff_1431
        assign out_data[1431] = lut_1431_out;
    end
    endgenerate
    
    
    
    // LUT : 1432
    wire [63:0] lut_1432_table = 64'b0000000000000000000000000000000000000000000000001011000010110001;
    wire [5:0] lut_1432_select = {
                             in_data[386],
                             in_data[276],
                             in_data[101],
                             in_data[296],
                             in_data[192],
                             in_data[552]};
    
    wire lut_1432_out = lut_1432_table[lut_1432_select];
    
    generate
    if ( USE_REG ) begin : ff_1432
        reg   lut_1432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1432_ff <= lut_1432_out;
            end
        end
        
        assign out_data[1432] = lut_1432_ff;
    end
    else begin : no_ff_1432
        assign out_data[1432] = lut_1432_out;
    end
    endgenerate
    
    
    
    // LUT : 1433
    wire [63:0] lut_1433_table = 64'b1111000001010000111100001111000011110100111101011111000111110101;
    wire [5:0] lut_1433_select = {
                             in_data[212],
                             in_data[710],
                             in_data[311],
                             in_data[315],
                             in_data[725],
                             in_data[593]};
    
    wire lut_1433_out = lut_1433_table[lut_1433_select];
    
    generate
    if ( USE_REG ) begin : ff_1433
        reg   lut_1433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1433_ff <= lut_1433_out;
            end
        end
        
        assign out_data[1433] = lut_1433_ff;
    end
    else begin : no_ff_1433
        assign out_data[1433] = lut_1433_out;
    end
    endgenerate
    
    
    
    // LUT : 1434
    wire [63:0] lut_1434_table = 64'b0101010101010101111100000101010101010101010101010101000001010101;
    wire [5:0] lut_1434_select = {
                             in_data[692],
                             in_data[102],
                             in_data[415],
                             in_data[484],
                             in_data[48],
                             in_data[376]};
    
    wire lut_1434_out = lut_1434_table[lut_1434_select];
    
    generate
    if ( USE_REG ) begin : ff_1434
        reg   lut_1434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1434_ff <= lut_1434_out;
            end
        end
        
        assign out_data[1434] = lut_1434_ff;
    end
    else begin : no_ff_1434
        assign out_data[1434] = lut_1434_out;
    end
    endgenerate
    
    
    
    // LUT : 1435
    wire [63:0] lut_1435_table = 64'b0000000000000000111100001111000011110000000000001111000011110000;
    wire [5:0] lut_1435_select = {
                             in_data[662],
                             in_data[524],
                             in_data[634],
                             in_data[457],
                             in_data[116],
                             in_data[617]};
    
    wire lut_1435_out = lut_1435_table[lut_1435_select];
    
    generate
    if ( USE_REG ) begin : ff_1435
        reg   lut_1435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1435_ff <= lut_1435_out;
            end
        end
        
        assign out_data[1435] = lut_1435_ff;
    end
    else begin : no_ff_1435
        assign out_data[1435] = lut_1435_out;
    end
    endgenerate
    
    
    
    // LUT : 1436
    wire [63:0] lut_1436_table = 64'b1101000000000000111100000100000011010000000000001111000000000000;
    wire [5:0] lut_1436_select = {
                             in_data[64],
                             in_data[249],
                             in_data[382],
                             in_data[211],
                             in_data[206],
                             in_data[57]};
    
    wire lut_1436_out = lut_1436_table[lut_1436_select];
    
    generate
    if ( USE_REG ) begin : ff_1436
        reg   lut_1436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1436_ff <= lut_1436_out;
            end
        end
        
        assign out_data[1436] = lut_1436_ff;
    end
    else begin : no_ff_1436
        assign out_data[1436] = lut_1436_out;
    end
    endgenerate
    
    
    
    // LUT : 1437
    wire [63:0] lut_1437_table = 64'b1111111111111010111111111111111111110000000000001111111111110000;
    wire [5:0] lut_1437_select = {
                             in_data[653],
                             in_data[436],
                             in_data[343],
                             in_data[456],
                             in_data[729],
                             in_data[514]};
    
    wire lut_1437_out = lut_1437_table[lut_1437_select];
    
    generate
    if ( USE_REG ) begin : ff_1437
        reg   lut_1437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1437_ff <= lut_1437_out;
            end
        end
        
        assign out_data[1437] = lut_1437_ff;
    end
    else begin : no_ff_1437
        assign out_data[1437] = lut_1437_out;
    end
    endgenerate
    
    
    
    // LUT : 1438
    wire [63:0] lut_1438_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_1438_select = {
                             in_data[339],
                             in_data[151],
                             in_data[548],
                             in_data[700],
                             in_data[19],
                             in_data[737]};
    
    wire lut_1438_out = lut_1438_table[lut_1438_select];
    
    generate
    if ( USE_REG ) begin : ff_1438
        reg   lut_1438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1438_ff <= lut_1438_out;
            end
        end
        
        assign out_data[1438] = lut_1438_ff;
    end
    else begin : no_ff_1438
        assign out_data[1438] = lut_1438_out;
    end
    endgenerate
    
    
    
    // LUT : 1439
    wire [63:0] lut_1439_table = 64'b1111111101010101111111111111111111001100010001000000100011001100;
    wire [5:0] lut_1439_select = {
                             in_data[323],
                             in_data[268],
                             in_data[539],
                             in_data[66],
                             in_data[220],
                             in_data[553]};
    
    wire lut_1439_out = lut_1439_table[lut_1439_select];
    
    generate
    if ( USE_REG ) begin : ff_1439
        reg   lut_1439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1439_ff <= lut_1439_out;
            end
        end
        
        assign out_data[1439] = lut_1439_ff;
    end
    else begin : no_ff_1439
        assign out_data[1439] = lut_1439_out;
    end
    endgenerate
    
    
    
    // LUT : 1440
    wire [63:0] lut_1440_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_1440_select = {
                             in_data[491],
                             in_data[696],
                             in_data[241],
                             in_data[767],
                             in_data[336],
                             in_data[559]};
    
    wire lut_1440_out = lut_1440_table[lut_1440_select];
    
    generate
    if ( USE_REG ) begin : ff_1440
        reg   lut_1440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1440_ff <= lut_1440_out;
            end
        end
        
        assign out_data[1440] = lut_1440_ff;
    end
    else begin : no_ff_1440
        assign out_data[1440] = lut_1440_out;
    end
    endgenerate
    
    
    
    // LUT : 1441
    wire [63:0] lut_1441_table = 64'b1111110111111101111111011111110111011000110111001101100011111100;
    wire [5:0] lut_1441_select = {
                             in_data[527],
                             in_data[252],
                             in_data[184],
                             in_data[164],
                             in_data[291],
                             in_data[495]};
    
    wire lut_1441_out = lut_1441_table[lut_1441_select];
    
    generate
    if ( USE_REG ) begin : ff_1441
        reg   lut_1441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1441_ff <= lut_1441_out;
            end
        end
        
        assign out_data[1441] = lut_1441_ff;
    end
    else begin : no_ff_1441
        assign out_data[1441] = lut_1441_out;
    end
    endgenerate
    
    
    
    // LUT : 1442
    wire [63:0] lut_1442_table = 64'b0100010011000100111111110100110101000100110001011100111111001101;
    wire [5:0] lut_1442_select = {
                             in_data[112],
                             in_data[349],
                             in_data[596],
                             in_data[213],
                             in_data[159],
                             in_data[682]};
    
    wire lut_1442_out = lut_1442_table[lut_1442_select];
    
    generate
    if ( USE_REG ) begin : ff_1442
        reg   lut_1442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1442_ff <= lut_1442_out;
            end
        end
        
        assign out_data[1442] = lut_1442_ff;
    end
    else begin : no_ff_1442
        assign out_data[1442] = lut_1442_out;
    end
    endgenerate
    
    
    
    // LUT : 1443
    wire [63:0] lut_1443_table = 64'b0000111000000000000000000000000011111111000000001111111100000000;
    wire [5:0] lut_1443_select = {
                             in_data[359],
                             in_data[592],
                             in_data[210],
                             in_data[367],
                             in_data[258],
                             in_data[21]};
    
    wire lut_1443_out = lut_1443_table[lut_1443_select];
    
    generate
    if ( USE_REG ) begin : ff_1443
        reg   lut_1443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1443_ff <= lut_1443_out;
            end
        end
        
        assign out_data[1443] = lut_1443_ff;
    end
    else begin : no_ff_1443
        assign out_data[1443] = lut_1443_out;
    end
    endgenerate
    
    
    
    // LUT : 1444
    wire [63:0] lut_1444_table = 64'b1111111111111111111111111111111100000000000000001011001010111010;
    wire [5:0] lut_1444_select = {
                             in_data[661],
                             in_data[607],
                             in_data[24],
                             in_data[74],
                             in_data[776],
                             in_data[158]};
    
    wire lut_1444_out = lut_1444_table[lut_1444_select];
    
    generate
    if ( USE_REG ) begin : ff_1444
        reg   lut_1444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1444_ff <= lut_1444_out;
            end
        end
        
        assign out_data[1444] = lut_1444_ff;
    end
    else begin : no_ff_1444
        assign out_data[1444] = lut_1444_out;
    end
    endgenerate
    
    
    
    // LUT : 1445
    wire [63:0] lut_1445_table = 64'b1111101111111111000000000000000010011001110111011000100011001000;
    wire [5:0] lut_1445_select = {
                             in_data[469],
                             in_data[432],
                             in_data[718],
                             in_data[389],
                             in_data[316],
                             in_data[594]};
    
    wire lut_1445_out = lut_1445_table[lut_1445_select];
    
    generate
    if ( USE_REG ) begin : ff_1445
        reg   lut_1445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1445_ff <= lut_1445_out;
            end
        end
        
        assign out_data[1445] = lut_1445_ff;
    end
    else begin : no_ff_1445
        assign out_data[1445] = lut_1445_out;
    end
    endgenerate
    
    
    
    // LUT : 1446
    wire [63:0] lut_1446_table = 64'b0000101000001010101010101010111100001010000010101010101010101011;
    wire [5:0] lut_1446_select = {
                             in_data[695],
                             in_data[269],
                             in_data[283],
                             in_data[465],
                             in_data[14],
                             in_data[602]};
    
    wire lut_1446_out = lut_1446_table[lut_1446_select];
    
    generate
    if ( USE_REG ) begin : ff_1446
        reg   lut_1446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1446_ff <= lut_1446_out;
            end
        end
        
        assign out_data[1446] = lut_1446_ff;
    end
    else begin : no_ff_1446
        assign out_data[1446] = lut_1446_out;
    end
    endgenerate
    
    
    
    // LUT : 1447
    wire [63:0] lut_1447_table = 64'b1000000010000000110111011101010110000000100000000101000111010001;
    wire [5:0] lut_1447_select = {
                             in_data[77],
                             in_data[470],
                             in_data[673],
                             in_data[375],
                             in_data[270],
                             in_data[581]};
    
    wire lut_1447_out = lut_1447_table[lut_1447_select];
    
    generate
    if ( USE_REG ) begin : ff_1447
        reg   lut_1447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1447_ff <= lut_1447_out;
            end
        end
        
        assign out_data[1447] = lut_1447_ff;
    end
    else begin : no_ff_1447
        assign out_data[1447] = lut_1447_out;
    end
    endgenerate
    
    
    
    // LUT : 1448
    wire [63:0] lut_1448_table = 64'b0010001000100010101110111011101000100010101010101011101011111110;
    wire [5:0] lut_1448_select = {
                             in_data[574],
                             in_data[288],
                             in_data[381],
                             in_data[32],
                             in_data[385],
                             in_data[629]};
    
    wire lut_1448_out = lut_1448_table[lut_1448_select];
    
    generate
    if ( USE_REG ) begin : ff_1448
        reg   lut_1448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1448_ff <= lut_1448_out;
            end
        end
        
        assign out_data[1448] = lut_1448_ff;
    end
    else begin : no_ff_1448
        assign out_data[1448] = lut_1448_out;
    end
    endgenerate
    
    
    
    // LUT : 1449
    wire [63:0] lut_1449_table = 64'b0001001100010011000100110001001100010011000100110001001100010011;
    wire [5:0] lut_1449_select = {
                             in_data[81],
                             in_data[39],
                             in_data[79],
                             in_data[666],
                             in_data[356],
                             in_data[409]};
    
    wire lut_1449_out = lut_1449_table[lut_1449_select];
    
    generate
    if ( USE_REG ) begin : ff_1449
        reg   lut_1449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1449_ff <= lut_1449_out;
            end
        end
        
        assign out_data[1449] = lut_1449_ff;
    end
    else begin : no_ff_1449
        assign out_data[1449] = lut_1449_out;
    end
    endgenerate
    
    
    
    // LUT : 1450
    wire [63:0] lut_1450_table = 64'b0111000111110101001100010111000101110001111101010011000101110001;
    wire [5:0] lut_1450_select = {
                             in_data[27],
                             in_data[750],
                             in_data[330],
                             in_data[719],
                             in_data[570],
                             in_data[471]};
    
    wire lut_1450_out = lut_1450_table[lut_1450_select];
    
    generate
    if ( USE_REG ) begin : ff_1450
        reg   lut_1450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1450_ff <= lut_1450_out;
            end
        end
        
        assign out_data[1450] = lut_1450_ff;
    end
    else begin : no_ff_1450
        assign out_data[1450] = lut_1450_out;
    end
    endgenerate
    
    
    
    // LUT : 1451
    wire [63:0] lut_1451_table = 64'b1010000000000000111100100000000011111111111111111111111111111111;
    wire [5:0] lut_1451_select = {
                             in_data[628],
                             in_data[165],
                             in_data[387],
                             in_data[468],
                             in_data[52],
                             in_data[34]};
    
    wire lut_1451_out = lut_1451_table[lut_1451_select];
    
    generate
    if ( USE_REG ) begin : ff_1451
        reg   lut_1451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1451_ff <= lut_1451_out;
            end
        end
        
        assign out_data[1451] = lut_1451_ff;
    end
    else begin : no_ff_1451
        assign out_data[1451] = lut_1451_out;
    end
    endgenerate
    
    
    
    // LUT : 1452
    wire [63:0] lut_1452_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1452_select = {
                             in_data[463],
                             in_data[772],
                             in_data[230],
                             in_data[11],
                             in_data[747],
                             in_data[257]};
    
    wire lut_1452_out = lut_1452_table[lut_1452_select];
    
    generate
    if ( USE_REG ) begin : ff_1452
        reg   lut_1452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1452_ff <= lut_1452_out;
            end
        end
        
        assign out_data[1452] = lut_1452_ff;
    end
    else begin : no_ff_1452
        assign out_data[1452] = lut_1452_out;
    end
    endgenerate
    
    
    
    // LUT : 1453
    wire [63:0] lut_1453_table = 64'b0000000000000000011101110111011100000000000000000111011101110111;
    wire [5:0] lut_1453_select = {
                             in_data[337],
                             in_data[413],
                             in_data[365],
                             in_data[616],
                             in_data[545],
                             in_data[649]};
    
    wire lut_1453_out = lut_1453_table[lut_1453_select];
    
    generate
    if ( USE_REG ) begin : ff_1453
        reg   lut_1453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1453_ff <= lut_1453_out;
            end
        end
        
        assign out_data[1453] = lut_1453_ff;
    end
    else begin : no_ff_1453
        assign out_data[1453] = lut_1453_out;
    end
    endgenerate
    
    
    
    // LUT : 1454
    wire [63:0] lut_1454_table = 64'b0000101011111111000000001111111010001010111111110000000011111110;
    wire [5:0] lut_1454_select = {
                             in_data[83],
                             in_data[485],
                             in_data[407],
                             in_data[410],
                             in_data[368],
                             in_data[603]};
    
    wire lut_1454_out = lut_1454_table[lut_1454_select];
    
    generate
    if ( USE_REG ) begin : ff_1454
        reg   lut_1454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1454_ff <= lut_1454_out;
            end
        end
        
        assign out_data[1454] = lut_1454_ff;
    end
    else begin : no_ff_1454
        assign out_data[1454] = lut_1454_out;
    end
    endgenerate
    
    
    
    // LUT : 1455
    wire [63:0] lut_1455_table = 64'b0000000000000000111111111111111100000000000000001111111111111111;
    wire [5:0] lut_1455_select = {
                             in_data[769],
                             in_data[515],
                             in_data[698],
                             in_data[50],
                             in_data[480],
                             in_data[782]};
    
    wire lut_1455_out = lut_1455_table[lut_1455_select];
    
    generate
    if ( USE_REG ) begin : ff_1455
        reg   lut_1455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1455_ff <= lut_1455_out;
            end
        end
        
        assign out_data[1455] = lut_1455_ff;
    end
    else begin : no_ff_1455
        assign out_data[1455] = lut_1455_out;
    end
    endgenerate
    
    
    
    // LUT : 1456
    wire [63:0] lut_1456_table = 64'b1000111011001110100010100000000011111111111111111110111111001100;
    wire [5:0] lut_1456_select = {
                             in_data[229],
                             in_data[711],
                             in_data[378],
                             in_data[199],
                             in_data[656],
                             in_data[218]};
    
    wire lut_1456_out = lut_1456_table[lut_1456_select];
    
    generate
    if ( USE_REG ) begin : ff_1456
        reg   lut_1456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1456_ff <= lut_1456_out;
            end
        end
        
        assign out_data[1456] = lut_1456_ff;
    end
    else begin : no_ff_1456
        assign out_data[1456] = lut_1456_out;
    end
    endgenerate
    
    
    
    // LUT : 1457
    wire [63:0] lut_1457_table = 64'b0000000000000000000000001110111100000000000000001111111111111111;
    wire [5:0] lut_1457_select = {
                             in_data[187],
                             in_data[156],
                             in_data[494],
                             in_data[78],
                             in_data[115],
                             in_data[306]};
    
    wire lut_1457_out = lut_1457_table[lut_1457_select];
    
    generate
    if ( USE_REG ) begin : ff_1457
        reg   lut_1457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1457_ff <= lut_1457_out;
            end
        end
        
        assign out_data[1457] = lut_1457_ff;
    end
    else begin : no_ff_1457
        assign out_data[1457] = lut_1457_out;
    end
    endgenerate
    
    
    
    // LUT : 1458
    wire [63:0] lut_1458_table = 64'b0011001111110011000000000010001000110011111100110000000000110010;
    wire [5:0] lut_1458_select = {
                             in_data[1],
                             in_data[430],
                             in_data[379],
                             in_data[106],
                             in_data[657],
                             in_data[780]};
    
    wire lut_1458_out = lut_1458_table[lut_1458_select];
    
    generate
    if ( USE_REG ) begin : ff_1458
        reg   lut_1458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1458_ff <= lut_1458_out;
            end
        end
        
        assign out_data[1458] = lut_1458_ff;
    end
    else begin : no_ff_1458
        assign out_data[1458] = lut_1458_out;
    end
    endgenerate
    
    
    
    // LUT : 1459
    wire [63:0] lut_1459_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1459_select = {
                             in_data[129],
                             in_data[401],
                             in_data[764],
                             in_data[771],
                             in_data[372],
                             in_data[614]};
    
    wire lut_1459_out = lut_1459_table[lut_1459_select];
    
    generate
    if ( USE_REG ) begin : ff_1459
        reg   lut_1459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1459_ff <= lut_1459_out;
            end
        end
        
        assign out_data[1459] = lut_1459_ff;
    end
    else begin : no_ff_1459
        assign out_data[1459] = lut_1459_out;
    end
    endgenerate
    
    
    
    // LUT : 1460
    wire [63:0] lut_1460_table = 64'b0000000000000000001010101010101000000000000000000010001010101010;
    wire [5:0] lut_1460_select = {
                             in_data[281],
                             in_data[554],
                             in_data[75],
                             in_data[86],
                             in_data[167],
                             in_data[461]};
    
    wire lut_1460_out = lut_1460_table[lut_1460_select];
    
    generate
    if ( USE_REG ) begin : ff_1460
        reg   lut_1460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1460_ff <= lut_1460_out;
            end
        end
        
        assign out_data[1460] = lut_1460_ff;
    end
    else begin : no_ff_1460
        assign out_data[1460] = lut_1460_out;
    end
    endgenerate
    
    
    
    // LUT : 1461
    wire [63:0] lut_1461_table = 64'b0000111100001111000011110000111100001101000011000000111100001111;
    wire [5:0] lut_1461_select = {
                             in_data[540],
                             in_data[76],
                             in_data[55],
                             in_data[209],
                             in_data[242],
                             in_data[777]};
    
    wire lut_1461_out = lut_1461_table[lut_1461_select];
    
    generate
    if ( USE_REG ) begin : ff_1461
        reg   lut_1461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1461_ff <= lut_1461_out;
            end
        end
        
        assign out_data[1461] = lut_1461_ff;
    end
    else begin : no_ff_1461
        assign out_data[1461] = lut_1461_out;
    end
    endgenerate
    
    
    
    // LUT : 1462
    wire [63:0] lut_1462_table = 64'b0101000001010000110101011101010011010100010100001111010111110101;
    wire [5:0] lut_1462_select = {
                             in_data[525],
                             in_data[131],
                             in_data[30],
                             in_data[295],
                             in_data[451],
                             in_data[486]};
    
    wire lut_1462_out = lut_1462_table[lut_1462_select];
    
    generate
    if ( USE_REG ) begin : ff_1462
        reg   lut_1462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1462_ff <= lut_1462_out;
            end
        end
        
        assign out_data[1462] = lut_1462_ff;
    end
    else begin : no_ff_1462
        assign out_data[1462] = lut_1462_out;
    end
    endgenerate
    
    
    
    // LUT : 1463
    wire [63:0] lut_1463_table = 64'b1111110011101100111111011111110111110100110100001111000001110001;
    wire [5:0] lut_1463_select = {
                             in_data[178],
                             in_data[260],
                             in_data[132],
                             in_data[526],
                             in_data[236],
                             in_data[689]};
    
    wire lut_1463_out = lut_1463_table[lut_1463_select];
    
    generate
    if ( USE_REG ) begin : ff_1463
        reg   lut_1463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1463_ff <= lut_1463_out;
            end
        end
        
        assign out_data[1463] = lut_1463_ff;
    end
    else begin : no_ff_1463
        assign out_data[1463] = lut_1463_out;
    end
    endgenerate
    
    
    
    // LUT : 1464
    wire [63:0] lut_1464_table = 64'b1010000010100000101010101011101011111010111110101111111111111011;
    wire [5:0] lut_1464_select = {
                             in_data[97],
                             in_data[194],
                             in_data[140],
                             in_data[109],
                             in_data[6],
                             in_data[650]};
    
    wire lut_1464_out = lut_1464_table[lut_1464_select];
    
    generate
    if ( USE_REG ) begin : ff_1464
        reg   lut_1464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1464_ff <= lut_1464_out;
            end
        end
        
        assign out_data[1464] = lut_1464_ff;
    end
    else begin : no_ff_1464
        assign out_data[1464] = lut_1464_out;
    end
    endgenerate
    
    
    
    // LUT : 1465
    wire [63:0] lut_1465_table = 64'b1010101101001101111111111101110100100010000000001000000000000000;
    wire [5:0] lut_1465_select = {
                             in_data[355],
                             in_data[152],
                             in_data[633],
                             in_data[473],
                             in_data[186],
                             in_data[541]};
    
    wire lut_1465_out = lut_1465_table[lut_1465_select];
    
    generate
    if ( USE_REG ) begin : ff_1465
        reg   lut_1465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1465_ff <= lut_1465_out;
            end
        end
        
        assign out_data[1465] = lut_1465_ff;
    end
    else begin : no_ff_1465
        assign out_data[1465] = lut_1465_out;
    end
    endgenerate
    
    
    
    // LUT : 1466
    wire [63:0] lut_1466_table = 64'b0000000000000000000000000000000000000000000000000101010101010101;
    wire [5:0] lut_1466_select = {
                             in_data[460],
                             in_data[93],
                             in_data[775],
                             in_data[779],
                             in_data[143],
                             in_data[191]};
    
    wire lut_1466_out = lut_1466_table[lut_1466_select];
    
    generate
    if ( USE_REG ) begin : ff_1466
        reg   lut_1466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1466_ff <= lut_1466_out;
            end
        end
        
        assign out_data[1466] = lut_1466_ff;
    end
    else begin : no_ff_1466
        assign out_data[1466] = lut_1466_out;
    end
    endgenerate
    
    
    
    // LUT : 1467
    wire [63:0] lut_1467_table = 64'b0111001111110001111111111111010101110001011100001111110111110100;
    wire [5:0] lut_1467_select = {
                             in_data[712],
                             in_data[153],
                             in_data[341],
                             in_data[176],
                             in_data[233],
                             in_data[161]};
    
    wire lut_1467_out = lut_1467_table[lut_1467_select];
    
    generate
    if ( USE_REG ) begin : ff_1467
        reg   lut_1467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1467_ff <= lut_1467_out;
            end
        end
        
        assign out_data[1467] = lut_1467_ff;
    end
    else begin : no_ff_1467
        assign out_data[1467] = lut_1467_out;
    end
    endgenerate
    
    
    
    // LUT : 1468
    wire [63:0] lut_1468_table = 64'b0000000000000000000000000000000011110101111101011111010111110100;
    wire [5:0] lut_1468_select = {
                             in_data[555],
                             in_data[25],
                             in_data[734],
                             in_data[183],
                             in_data[100],
                             in_data[572]};
    
    wire lut_1468_out = lut_1468_table[lut_1468_select];
    
    generate
    if ( USE_REG ) begin : ff_1468
        reg   lut_1468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1468_ff <= lut_1468_out;
            end
        end
        
        assign out_data[1468] = lut_1468_ff;
    end
    else begin : no_ff_1468
        assign out_data[1468] = lut_1468_out;
    end
    endgenerate
    
    
    
    // LUT : 1469
    wire [63:0] lut_1469_table = 64'b0000000000000000010101010101010100000000000000001111010111110101;
    wire [5:0] lut_1469_select = {
                             in_data[207],
                             in_data[637],
                             in_data[362],
                             in_data[340],
                             in_data[450],
                             in_data[605]};
    
    wire lut_1469_out = lut_1469_table[lut_1469_select];
    
    generate
    if ( USE_REG ) begin : ff_1469
        reg   lut_1469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1469_ff <= lut_1469_out;
            end
        end
        
        assign out_data[1469] = lut_1469_ff;
    end
    else begin : no_ff_1469
        assign out_data[1469] = lut_1469_out;
    end
    endgenerate
    
    
    
    // LUT : 1470
    wire [63:0] lut_1470_table = 64'b0000001100001011000000110000101100001011000010110000101100001111;
    wire [5:0] lut_1470_select = {
                             in_data[88],
                             in_data[762],
                             in_data[40],
                             in_data[431],
                             in_data[265],
                             in_data[697]};
    
    wire lut_1470_out = lut_1470_table[lut_1470_select];
    
    generate
    if ( USE_REG ) begin : ff_1470
        reg   lut_1470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1470_ff <= lut_1470_out;
            end
        end
        
        assign out_data[1470] = lut_1470_ff;
    end
    else begin : no_ff_1470
        assign out_data[1470] = lut_1470_out;
    end
    endgenerate
    
    
    
    // LUT : 1471
    wire [63:0] lut_1471_table = 64'b1111011111110111111100011111000111110111111101111111000111110001;
    wire [5:0] lut_1471_select = {
                             in_data[781],
                             in_data[678],
                             in_data[643],
                             in_data[174],
                             in_data[403],
                             in_data[440]};
    
    wire lut_1471_out = lut_1471_table[lut_1471_select];
    
    generate
    if ( USE_REG ) begin : ff_1471
        reg   lut_1471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1471_ff <= lut_1471_out;
            end
        end
        
        assign out_data[1471] = lut_1471_ff;
    end
    else begin : no_ff_1471
        assign out_data[1471] = lut_1471_out;
    end
    endgenerate
    
    
    
    // LUT : 1472
    wire [63:0] lut_1472_table = 64'b1110111011101110111010001110100011111111111111111111111111111111;
    wire [5:0] lut_1472_select = {
                             in_data[380],
                             in_data[371],
                             in_data[13],
                             in_data[738],
                             in_data[556],
                             in_data[648]};
    
    wire lut_1472_out = lut_1472_table[lut_1472_select];
    
    generate
    if ( USE_REG ) begin : ff_1472
        reg   lut_1472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1472_ff <= lut_1472_out;
            end
        end
        
        assign out_data[1472] = lut_1472_ff;
    end
    else begin : no_ff_1472
        assign out_data[1472] = lut_1472_out;
    end
    endgenerate
    
    
    
    // LUT : 1473
    wire [63:0] lut_1473_table = 64'b0000000000000000000100010101000100000000000000000111010111110111;
    wire [5:0] lut_1473_select = {
                             in_data[479],
                             in_data[437],
                             in_data[704],
                             in_data[369],
                             in_data[266],
                             in_data[550]};
    
    wire lut_1473_out = lut_1473_table[lut_1473_select];
    
    generate
    if ( USE_REG ) begin : ff_1473
        reg   lut_1473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1473_ff <= lut_1473_out;
            end
        end
        
        assign out_data[1473] = lut_1473_ff;
    end
    else begin : no_ff_1473
        assign out_data[1473] = lut_1473_out;
    end
    endgenerate
    
    
    
    // LUT : 1474
    wire [63:0] lut_1474_table = 64'b1010101010101010111111111111111110101010101010101111111111111111;
    wire [5:0] lut_1474_select = {
                             in_data[417],
                             in_data[571],
                             in_data[641],
                             in_data[744],
                             in_data[363],
                             in_data[424]};
    
    wire lut_1474_out = lut_1474_table[lut_1474_select];
    
    generate
    if ( USE_REG ) begin : ff_1474
        reg   lut_1474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1474_ff <= lut_1474_out;
            end
        end
        
        assign out_data[1474] = lut_1474_ff;
    end
    else begin : no_ff_1474
        assign out_data[1474] = lut_1474_out;
    end
    endgenerate
    
    
    
    // LUT : 1475
    wire [63:0] lut_1475_table = 64'b0000000000000000000000000000000011100000111111101110000011111110;
    wire [5:0] lut_1475_select = {
                             in_data[294],
                             in_data[560],
                             in_data[624],
                             in_data[263],
                             in_data[72],
                             in_data[397]};
    
    wire lut_1475_out = lut_1475_table[lut_1475_select];
    
    generate
    if ( USE_REG ) begin : ff_1475
        reg   lut_1475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1475_ff <= lut_1475_out;
            end
        end
        
        assign out_data[1475] = lut_1475_ff;
    end
    else begin : no_ff_1475
        assign out_data[1475] = lut_1475_out;
    end
    endgenerate
    
    
    
    // LUT : 1476
    wire [63:0] lut_1476_table = 64'b0000000000100000111110111111101100000000000000001011001111110011;
    wire [5:0] lut_1476_select = {
                             in_data[227],
                             in_data[582],
                             in_data[390],
                             in_data[622],
                             in_data[318],
                             in_data[478]};
    
    wire lut_1476_out = lut_1476_table[lut_1476_select];
    
    generate
    if ( USE_REG ) begin : ff_1476
        reg   lut_1476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1476_ff <= lut_1476_out;
            end
        end
        
        assign out_data[1476] = lut_1476_ff;
    end
    else begin : no_ff_1476
        assign out_data[1476] = lut_1476_out;
    end
    endgenerate
    
    
    
    // LUT : 1477
    wire [63:0] lut_1477_table = 64'b0011000100110001110100001101000000110011001100111111000011010100;
    wire [5:0] lut_1477_select = {
                             in_data[248],
                             in_data[499],
                             in_data[23],
                             in_data[496],
                             in_data[352],
                             in_data[577]};
    
    wire lut_1477_out = lut_1477_table[lut_1477_select];
    
    generate
    if ( USE_REG ) begin : ff_1477
        reg   lut_1477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1477_ff <= lut_1477_out;
            end
        end
        
        assign out_data[1477] = lut_1477_ff;
    end
    else begin : no_ff_1477
        assign out_data[1477] = lut_1477_out;
    end
    endgenerate
    
    
    
    // LUT : 1478
    wire [63:0] lut_1478_table = 64'b1111111100000000111111110000000011110001000000001111001100000000;
    wire [5:0] lut_1478_select = {
                             in_data[217],
                             in_data[590],
                             in_data[489],
                             in_data[685],
                             in_data[620],
                             in_data[416]};
    
    wire lut_1478_out = lut_1478_table[lut_1478_select];
    
    generate
    if ( USE_REG ) begin : ff_1478
        reg   lut_1478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1478_ff <= lut_1478_out;
            end
        end
        
        assign out_data[1478] = lut_1478_ff;
    end
    else begin : no_ff_1478
        assign out_data[1478] = lut_1478_out;
    end
    endgenerate
    
    
    
    // LUT : 1479
    wire [63:0] lut_1479_table = 64'b0000000011111111000000001111111111101111111111110000000000001111;
    wire [5:0] lut_1479_select = {
                             in_data[488],
                             in_data[442],
                             in_data[235],
                             in_data[395],
                             in_data[504],
                             in_data[671]};
    
    wire lut_1479_out = lut_1479_table[lut_1479_select];
    
    generate
    if ( USE_REG ) begin : ff_1479
        reg   lut_1479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1479_ff <= lut_1479_out;
            end
        end
        
        assign out_data[1479] = lut_1479_ff;
    end
    else begin : no_ff_1479
        assign out_data[1479] = lut_1479_out;
    end
    endgenerate
    
    
    
    // LUT : 1480
    wire [63:0] lut_1480_table = 64'b1111111111111111101010101010101011111111111111111010101010101010;
    wire [5:0] lut_1480_select = {
                             in_data[225],
                             in_data[103],
                             in_data[783],
                             in_data[672],
                             in_data[334],
                             in_data[154]};
    
    wire lut_1480_out = lut_1480_table[lut_1480_select];
    
    generate
    if ( USE_REG ) begin : ff_1480
        reg   lut_1480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1480_ff <= lut_1480_out;
            end
        end
        
        assign out_data[1480] = lut_1480_ff;
    end
    else begin : no_ff_1480
        assign out_data[1480] = lut_1480_out;
    end
    endgenerate
    
    
    
    // LUT : 1481
    wire [63:0] lut_1481_table = 64'b0000000000000000111100001111001100000000000000001111000011110000;
    wire [5:0] lut_1481_select = {
                             in_data[46],
                             in_data[68],
                             in_data[90],
                             in_data[180],
                             in_data[166],
                             in_data[92]};
    
    wire lut_1481_out = lut_1481_table[lut_1481_select];
    
    generate
    if ( USE_REG ) begin : ff_1481
        reg   lut_1481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1481_ff <= lut_1481_out;
            end
        end
        
        assign out_data[1481] = lut_1481_ff;
    end
    else begin : no_ff_1481
        assign out_data[1481] = lut_1481_out;
    end
    endgenerate
    
    
    
    // LUT : 1482
    wire [63:0] lut_1482_table = 64'b1111101111111010111110101111101011110010111110101111001011111010;
    wire [5:0] lut_1482_select = {
                             in_data[214],
                             in_data[575],
                             in_data[182],
                             in_data[568],
                             in_data[261],
                             in_data[127]};
    
    wire lut_1482_out = lut_1482_table[lut_1482_select];
    
    generate
    if ( USE_REG ) begin : ff_1482
        reg   lut_1482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1482_ff <= lut_1482_out;
            end
        end
        
        assign out_data[1482] = lut_1482_ff;
    end
    else begin : no_ff_1482
        assign out_data[1482] = lut_1482_out;
    end
    endgenerate
    
    
    
    // LUT : 1483
    wire [63:0] lut_1483_table = 64'b1111100011111000111110001111100011111000111110001111100011111000;
    wire [5:0] lut_1483_select = {
                             in_data[752],
                             in_data[224],
                             in_data[758],
                             in_data[322],
                             in_data[635],
                             in_data[344]};
    
    wire lut_1483_out = lut_1483_table[lut_1483_select];
    
    generate
    if ( USE_REG ) begin : ff_1483
        reg   lut_1483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1483_ff <= lut_1483_out;
            end
        end
        
        assign out_data[1483] = lut_1483_ff;
    end
    else begin : no_ff_1483
        assign out_data[1483] = lut_1483_out;
    end
    endgenerate
    
    
    
    // LUT : 1484
    wire [63:0] lut_1484_table = 64'b0000010011001100000001001100110000000000010001010000010101010101;
    wire [5:0] lut_1484_select = {
                             in_data[467],
                             in_data[41],
                             in_data[126],
                             in_data[284],
                             in_data[472],
                             in_data[208]};
    
    wire lut_1484_out = lut_1484_table[lut_1484_select];
    
    generate
    if ( USE_REG ) begin : ff_1484
        reg   lut_1484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1484_ff <= lut_1484_out;
            end
        end
        
        assign out_data[1484] = lut_1484_ff;
    end
    else begin : no_ff_1484
        assign out_data[1484] = lut_1484_out;
    end
    endgenerate
    
    
    
    // LUT : 1485
    wire [63:0] lut_1485_table = 64'b0000000000000000000000000000000011111111111111111111001011111011;
    wire [5:0] lut_1485_select = {
                             in_data[320],
                             in_data[117],
                             in_data[85],
                             in_data[353],
                             in_data[354],
                             in_data[392]};
    
    wire lut_1485_out = lut_1485_table[lut_1485_select];
    
    generate
    if ( USE_REG ) begin : ff_1485
        reg   lut_1485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1485_ff <= lut_1485_out;
            end
        end
        
        assign out_data[1485] = lut_1485_ff;
    end
    else begin : no_ff_1485
        assign out_data[1485] = lut_1485_out;
    end
    endgenerate
    
    
    
    // LUT : 1486
    wire [63:0] lut_1486_table = 64'b0000000000000000000000000101010100000000000000000000000101010101;
    wire [5:0] lut_1486_select = {
                             in_data[538],
                             in_data[452],
                             in_data[474],
                             in_data[705],
                             in_data[80],
                             in_data[243]};
    
    wire lut_1486_out = lut_1486_table[lut_1486_select];
    
    generate
    if ( USE_REG ) begin : ff_1486
        reg   lut_1486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1486_ff <= lut_1486_out;
            end
        end
        
        assign out_data[1486] = lut_1486_ff;
    end
    else begin : no_ff_1486
        assign out_data[1486] = lut_1486_out;
    end
    endgenerate
    
    
    
    // LUT : 1487
    wire [63:0] lut_1487_table = 64'b0000000000000000000010100000000000001010000000001111111101011111;
    wire [5:0] lut_1487_select = {
                             in_data[221],
                             in_data[350],
                             in_data[324],
                             in_data[523],
                             in_data[675],
                             in_data[237]};
    
    wire lut_1487_out = lut_1487_table[lut_1487_select];
    
    generate
    if ( USE_REG ) begin : ff_1487
        reg   lut_1487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1487_ff <= lut_1487_out;
            end
        end
        
        assign out_data[1487] = lut_1487_ff;
    end
    else begin : no_ff_1487
        assign out_data[1487] = lut_1487_out;
    end
    endgenerate
    
    
    
    // LUT : 1488
    wire [63:0] lut_1488_table = 64'b1111111111111111111111111111111111111111111111111010101010101010;
    wire [5:0] lut_1488_select = {
                             in_data[128],
                             in_data[683],
                             in_data[63],
                             in_data[84],
                             in_data[169],
                             in_data[44]};
    
    wire lut_1488_out = lut_1488_table[lut_1488_select];
    
    generate
    if ( USE_REG ) begin : ff_1488
        reg   lut_1488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1488_ff <= lut_1488_out;
            end
        end
        
        assign out_data[1488] = lut_1488_ff;
    end
    else begin : no_ff_1488
        assign out_data[1488] = lut_1488_out;
    end
    endgenerate
    
    
    
    // LUT : 1489
    wire [63:0] lut_1489_table = 64'b0101010011111111010101011111111101000100110111110100010011011101;
    wire [5:0] lut_1489_select = {
                             in_data[297],
                             in_data[561],
                             in_data[408],
                             in_data[60],
                             in_data[203],
                             in_data[722]};
    
    wire lut_1489_out = lut_1489_table[lut_1489_select];
    
    generate
    if ( USE_REG ) begin : ff_1489
        reg   lut_1489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1489_ff <= lut_1489_out;
            end
        end
        
        assign out_data[1489] = lut_1489_ff;
    end
    else begin : no_ff_1489
        assign out_data[1489] = lut_1489_out;
    end
    endgenerate
    
    
    
    // LUT : 1490
    wire [63:0] lut_1490_table = 64'b0000000001010000000000000010000001010000010100000000000001010000;
    wire [5:0] lut_1490_select = {
                             in_data[597],
                             in_data[314],
                             in_data[501],
                             in_data[466],
                             in_data[608],
                             in_data[598]};
    
    wire lut_1490_out = lut_1490_table[lut_1490_select];
    
    generate
    if ( USE_REG ) begin : ff_1490
        reg   lut_1490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1490_ff <= lut_1490_out;
            end
        end
        
        assign out_data[1490] = lut_1490_ff;
    end
    else begin : no_ff_1490
        assign out_data[1490] = lut_1490_out;
    end
    endgenerate
    
    
    
    // LUT : 1491
    wire [63:0] lut_1491_table = 64'b0011001111111011001100111111101100000011000000110000001100000011;
    wire [5:0] lut_1491_select = {
                             in_data[175],
                             in_data[308],
                             in_data[134],
                             in_data[238],
                             in_data[373],
                             in_data[37]};
    
    wire lut_1491_out = lut_1491_table[lut_1491_select];
    
    generate
    if ( USE_REG ) begin : ff_1491
        reg   lut_1491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1491_ff <= lut_1491_out;
            end
        end
        
        assign out_data[1491] = lut_1491_ff;
    end
    else begin : no_ff_1491
        assign out_data[1491] = lut_1491_out;
    end
    endgenerate
    
    
    
    // LUT : 1492
    wire [63:0] lut_1492_table = 64'b1111111111001100000000000100010111011101110011000000000011001101;
    wire [5:0] lut_1492_select = {
                             in_data[500],
                             in_data[438],
                             in_data[406],
                             in_data[35],
                             in_data[516],
                             in_data[388]};
    
    wire lut_1492_out = lut_1492_table[lut_1492_select];
    
    generate
    if ( USE_REG ) begin : ff_1492
        reg   lut_1492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1492_ff <= lut_1492_out;
            end
        end
        
        assign out_data[1492] = lut_1492_ff;
    end
    else begin : no_ff_1492
        assign out_data[1492] = lut_1492_out;
    end
    endgenerate
    
    
    
    // LUT : 1493
    wire [63:0] lut_1493_table = 64'b1111111110111111111111111011101111111111101110111111111110111011;
    wire [5:0] lut_1493_select = {
                             in_data[82],
                             in_data[611],
                             in_data[148],
                             in_data[348],
                             in_data[383],
                             in_data[536]};
    
    wire lut_1493_out = lut_1493_table[lut_1493_select];
    
    generate
    if ( USE_REG ) begin : ff_1493
        reg   lut_1493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1493_ff <= lut_1493_out;
            end
        end
        
        assign out_data[1493] = lut_1493_ff;
    end
    else begin : no_ff_1493
        assign out_data[1493] = lut_1493_out;
    end
    endgenerate
    
    
    
    // LUT : 1494
    wire [63:0] lut_1494_table = 64'b0000000001010111000000000000000000000000111111111111111100000001;
    wire [5:0] lut_1494_select = {
                             in_data[275],
                             in_data[231],
                             in_data[609],
                             in_data[419],
                             in_data[732],
                             in_data[454]};
    
    wire lut_1494_out = lut_1494_table[lut_1494_select];
    
    generate
    if ( USE_REG ) begin : ff_1494
        reg   lut_1494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1494_ff <= lut_1494_out;
            end
        end
        
        assign out_data[1494] = lut_1494_ff;
    end
    else begin : no_ff_1494
        assign out_data[1494] = lut_1494_out;
    end
    endgenerate
    
    
    
    // LUT : 1495
    wire [63:0] lut_1495_table = 64'b0000000000000101000000000000000100000000000000000000000000000001;
    wire [5:0] lut_1495_select = {
                             in_data[721],
                             in_data[422],
                             in_data[667],
                             in_data[418],
                             in_data[585],
                             in_data[122]};
    
    wire lut_1495_out = lut_1495_table[lut_1495_select];
    
    generate
    if ( USE_REG ) begin : ff_1495
        reg   lut_1495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1495_ff <= lut_1495_out;
            end
        end
        
        assign out_data[1495] = lut_1495_ff;
    end
    else begin : no_ff_1495
        assign out_data[1495] = lut_1495_out;
    end
    endgenerate
    
    
    
    // LUT : 1496
    wire [63:0] lut_1496_table = 64'b1111111100001111000000000000000000001111000011110000000000000101;
    wire [5:0] lut_1496_select = {
                             in_data[293],
                             in_data[244],
                             in_data[483],
                             in_data[481],
                             in_data[0],
                             in_data[145]};
    
    wire lut_1496_out = lut_1496_table[lut_1496_select];
    
    generate
    if ( USE_REG ) begin : ff_1496
        reg   lut_1496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1496_ff <= lut_1496_out;
            end
        end
        
        assign out_data[1496] = lut_1496_ff;
    end
    else begin : no_ff_1496
        assign out_data[1496] = lut_1496_out;
    end
    endgenerate
    
    
    
    // LUT : 1497
    wire [63:0] lut_1497_table = 64'b0111011100110011010111110011001111111100111111111111110011111111;
    wire [5:0] lut_1497_select = {
                             in_data[549],
                             in_data[476],
                             in_data[517],
                             in_data[565],
                             in_data[604],
                             in_data[551]};
    
    wire lut_1497_out = lut_1497_table[lut_1497_select];
    
    generate
    if ( USE_REG ) begin : ff_1497
        reg   lut_1497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1497_ff <= lut_1497_out;
            end
        end
        
        assign out_data[1497] = lut_1497_ff;
    end
    else begin : no_ff_1497
        assign out_data[1497] = lut_1497_out;
    end
    endgenerate
    
    
    
    // LUT : 1498
    wire [63:0] lut_1498_table = 64'b0000000000000101111100001111000000000000000001011111000011110000;
    wire [5:0] lut_1498_select = {
                             in_data[53],
                             in_data[292],
                             in_data[247],
                             in_data[271],
                             in_data[642],
                             in_data[591]};
    
    wire lut_1498_out = lut_1498_table[lut_1498_select];
    
    generate
    if ( USE_REG ) begin : ff_1498
        reg   lut_1498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1498_ff <= lut_1498_out;
            end
        end
        
        assign out_data[1498] = lut_1498_ff;
    end
    else begin : no_ff_1498
        assign out_data[1498] = lut_1498_out;
    end
    endgenerate
    
    
    
    // LUT : 1499
    wire [63:0] lut_1499_table = 64'b1010000011101000101010101111111110101010111010101111111011111111;
    wire [5:0] lut_1499_select = {
                             in_data[428],
                             in_data[347],
                             in_data[185],
                             in_data[706],
                             in_data[576],
                             in_data[299]};
    
    wire lut_1499_out = lut_1499_table[lut_1499_select];
    
    generate
    if ( USE_REG ) begin : ff_1499
        reg   lut_1499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1499_ff <= lut_1499_out;
            end
        end
        
        assign out_data[1499] = lut_1499_ff;
    end
    else begin : no_ff_1499
        assign out_data[1499] = lut_1499_out;
    end
    endgenerate
    
    
    
    // LUT : 1500
    wire [63:0] lut_1500_table = 64'b0000000000001111000000000010111100000000000011110000000000001111;
    wire [5:0] lut_1500_select = {
                             in_data[20],
                             in_data[364],
                             in_data[272],
                             in_data[250],
                             in_data[58],
                             in_data[507]};
    
    wire lut_1500_out = lut_1500_table[lut_1500_select];
    
    generate
    if ( USE_REG ) begin : ff_1500
        reg   lut_1500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1500_ff <= lut_1500_out;
            end
        end
        
        assign out_data[1500] = lut_1500_ff;
    end
    else begin : no_ff_1500
        assign out_data[1500] = lut_1500_out;
    end
    endgenerate
    
    
    
    // LUT : 1501
    wire [63:0] lut_1501_table = 64'b0000000000000011000000000000001100000000000000110000000000000011;
    wire [5:0] lut_1501_select = {
                             in_data[759],
                             in_data[669],
                             in_data[601],
                             in_data[528],
                             in_data[557],
                             in_data[703]};
    
    wire lut_1501_out = lut_1501_table[lut_1501_select];
    
    generate
    if ( USE_REG ) begin : ff_1501
        reg   lut_1501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1501_ff <= lut_1501_out;
            end
        end
        
        assign out_data[1501] = lut_1501_ff;
    end
    else begin : no_ff_1501
        assign out_data[1501] = lut_1501_out;
    end
    endgenerate
    
    
    
    // LUT : 1502
    wire [63:0] lut_1502_table = 64'b1111111111111111111111111111111100000000000000001101010011110100;
    wire [5:0] lut_1502_select = {
                             in_data[623],
                             in_data[190],
                             in_data[701],
                             in_data[120],
                             in_data[446],
                             in_data[709]};
    
    wire lut_1502_out = lut_1502_table[lut_1502_select];
    
    generate
    if ( USE_REG ) begin : ff_1502
        reg   lut_1502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1502_ff <= lut_1502_out;
            end
        end
        
        assign out_data[1502] = lut_1502_ff;
    end
    else begin : no_ff_1502
        assign out_data[1502] = lut_1502_out;
    end
    endgenerate
    
    
    
    // LUT : 1503
    wire [63:0] lut_1503_table = 64'b1010000011101000111000001110100011101110111011101110111011101111;
    wire [5:0] lut_1503_select = {
                             in_data[179],
                             in_data[61],
                             in_data[563],
                             in_data[578],
                             in_data[482],
                             in_data[313]};
    
    wire lut_1503_out = lut_1503_table[lut_1503_select];
    
    generate
    if ( USE_REG ) begin : ff_1503
        reg   lut_1503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1503_ff <= lut_1503_out;
            end
        end
        
        assign out_data[1503] = lut_1503_ff;
    end
    else begin : no_ff_1503
        assign out_data[1503] = lut_1503_out;
    end
    endgenerate
    
    
    
    // LUT : 1504
    wire [63:0] lut_1504_table = 64'b0000000000000000000000000000000000000000000000000101010101010101;
    wire [5:0] lut_1504_select = {
                             in_data[498],
                             in_data[691],
                             in_data[28],
                             in_data[312],
                             in_data[778],
                             in_data[717]};
    
    wire lut_1504_out = lut_1504_table[lut_1504_select];
    
    generate
    if ( USE_REG ) begin : ff_1504
        reg   lut_1504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1504_ff <= lut_1504_out;
            end
        end
        
        assign out_data[1504] = lut_1504_ff;
    end
    else begin : no_ff_1504
        assign out_data[1504] = lut_1504_out;
    end
    endgenerate
    
    
    
    // LUT : 1505
    wire [63:0] lut_1505_table = 64'b0000000000000000000000000000000001111111010101010101010101010101;
    wire [5:0] lut_1505_select = {
                             in_data[606],
                             in_data[22],
                             in_data[319],
                             in_data[421],
                             in_data[646],
                             in_data[123]};
    
    wire lut_1505_out = lut_1505_table[lut_1505_select];
    
    generate
    if ( USE_REG ) begin : ff_1505
        reg   lut_1505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1505_ff <= lut_1505_out;
            end
        end
        
        assign out_data[1505] = lut_1505_ff;
    end
    else begin : no_ff_1505
        assign out_data[1505] = lut_1505_out;
    end
    endgenerate
    
    
    
    // LUT : 1506
    wire [63:0] lut_1506_table = 64'b1111001111111111111000001111110011110011111111111110000011111000;
    wire [5:0] lut_1506_select = {
                             in_data[588],
                             in_data[267],
                             in_data[716],
                             in_data[118],
                             in_data[537],
                             in_data[612]};
    
    wire lut_1506_out = lut_1506_table[lut_1506_select];
    
    generate
    if ( USE_REG ) begin : ff_1506
        reg   lut_1506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1506_ff <= lut_1506_out;
            end
        end
        
        assign out_data[1506] = lut_1506_ff;
    end
    else begin : no_ff_1506
        assign out_data[1506] = lut_1506_out;
    end
    endgenerate
    
    
    
    // LUT : 1507
    wire [63:0] lut_1507_table = 64'b0000000001110011000000000111001100000000001100110000000000111011;
    wire [5:0] lut_1507_select = {
                             in_data[5],
                             in_data[279],
                             in_data[99],
                             in_data[645],
                             in_data[400],
                             in_data[168]};
    
    wire lut_1507_out = lut_1507_table[lut_1507_select];
    
    generate
    if ( USE_REG ) begin : ff_1507
        reg   lut_1507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1507_ff <= lut_1507_out;
            end
        end
        
        assign out_data[1507] = lut_1507_ff;
    end
    else begin : no_ff_1507
        assign out_data[1507] = lut_1507_out;
    end
    endgenerate
    
    
    
    // LUT : 1508
    wire [63:0] lut_1508_table = 64'b1111111111111111010100000001000011111111111111110001000000010000;
    wire [5:0] lut_1508_select = {
                             in_data[615],
                             in_data[511],
                             in_data[477],
                             in_data[326],
                             in_data[73],
                             in_data[506]};
    
    wire lut_1508_out = lut_1508_table[lut_1508_select];
    
    generate
    if ( USE_REG ) begin : ff_1508
        reg   lut_1508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1508_ff <= lut_1508_out;
            end
        end
        
        assign out_data[1508] = lut_1508_ff;
    end
    else begin : no_ff_1508
        assign out_data[1508] = lut_1508_out;
    end
    endgenerate
    
    
    
    // LUT : 1509
    wire [63:0] lut_1509_table = 64'b1110111111101111111111111111111100000000000010001000100010000000;
    wire [5:0] lut_1509_select = {
                             in_data[439],
                             in_data[105],
                             in_data[36],
                             in_data[160],
                             in_data[228],
                             in_data[232]};
    
    wire lut_1509_out = lut_1509_table[lut_1509_select];
    
    generate
    if ( USE_REG ) begin : ff_1509
        reg   lut_1509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1509_ff <= lut_1509_out;
            end
        end
        
        assign out_data[1509] = lut_1509_ff;
    end
    else begin : no_ff_1509
        assign out_data[1509] = lut_1509_out;
    end
    endgenerate
    
    
    
    // LUT : 1510
    wire [63:0] lut_1510_table = 64'b0101010100010000010101010101000000000101000000000101010100010101;
    wire [5:0] lut_1510_select = {
                             in_data[287],
                             in_data[509],
                             in_data[544],
                             in_data[119],
                             in_data[18],
                             in_data[659]};
    
    wire lut_1510_out = lut_1510_table[lut_1510_select];
    
    generate
    if ( USE_REG ) begin : ff_1510
        reg   lut_1510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1510_ff <= lut_1510_out;
            end
        end
        
        assign out_data[1510] = lut_1510_ff;
    end
    else begin : no_ff_1510
        assign out_data[1510] = lut_1510_out;
    end
    endgenerate
    
    
    
    // LUT : 1511
    wire [63:0] lut_1511_table = 64'b1111111111111111000000000000000011111111111111110000101100001010;
    wire [5:0] lut_1511_select = {
                             in_data[462],
                             in_data[411],
                             in_data[7],
                             in_data[619],
                             in_data[195],
                             in_data[763]};
    
    wire lut_1511_out = lut_1511_table[lut_1511_select];
    
    generate
    if ( USE_REG ) begin : ff_1511
        reg   lut_1511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1511_ff <= lut_1511_out;
            end
        end
        
        assign out_data[1511] = lut_1511_ff;
    end
    else begin : no_ff_1511
        assign out_data[1511] = lut_1511_out;
    end
    endgenerate
    
    
    
    // LUT : 1512
    wire [63:0] lut_1512_table = 64'b1100110011001111110011001100111011001100110011111100110011001100;
    wire [5:0] lut_1512_select = {
                             in_data[532],
                             in_data[331],
                             in_data[425],
                             in_data[529],
                             in_data[681],
                             in_data[505]};
    
    wire lut_1512_out = lut_1512_table[lut_1512_select];
    
    generate
    if ( USE_REG ) begin : ff_1512
        reg   lut_1512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1512_ff <= lut_1512_out;
            end
        end
        
        assign out_data[1512] = lut_1512_ff;
    end
    else begin : no_ff_1512
        assign out_data[1512] = lut_1512_out;
    end
    endgenerate
    
    
    
    // LUT : 1513
    wire [63:0] lut_1513_table = 64'b0001000000010000000100000001000000010000000100010001000000010001;
    wire [5:0] lut_1513_select = {
                             in_data[731],
                             in_data[54],
                             in_data[307],
                             in_data[137],
                             in_data[742],
                             in_data[226]};
    
    wire lut_1513_out = lut_1513_table[lut_1513_select];
    
    generate
    if ( USE_REG ) begin : ff_1513
        reg   lut_1513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1513_ff <= lut_1513_out;
            end
        end
        
        assign out_data[1513] = lut_1513_ff;
    end
    else begin : no_ff_1513
        assign out_data[1513] = lut_1513_out;
    end
    endgenerate
    
    
    
    // LUT : 1514
    wire [63:0] lut_1514_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_1514_select = {
                             in_data[434],
                             in_data[328],
                             in_data[765],
                             in_data[8],
                             in_data[558],
                             in_data[332]};
    
    wire lut_1514_out = lut_1514_table[lut_1514_select];
    
    generate
    if ( USE_REG ) begin : ff_1514
        reg   lut_1514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1514_ff <= lut_1514_out;
            end
        end
        
        assign out_data[1514] = lut_1514_ff;
    end
    else begin : no_ff_1514
        assign out_data[1514] = lut_1514_out;
    end
    endgenerate
    
    
    
    // LUT : 1515
    wire [63:0] lut_1515_table = 64'b1111111100000000111111110000001111111111000000001111111100000011;
    wire [5:0] lut_1515_select = {
                             in_data[62],
                             in_data[453],
                             in_data[567],
                             in_data[610],
                             in_data[300],
                             in_data[33]};
    
    wire lut_1515_out = lut_1515_table[lut_1515_select];
    
    generate
    if ( USE_REG ) begin : ff_1515
        reg   lut_1515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1515_ff <= lut_1515_out;
            end
        end
        
        assign out_data[1515] = lut_1515_ff;
    end
    else begin : no_ff_1515
        assign out_data[1515] = lut_1515_out;
    end
    endgenerate
    
    
    
    // LUT : 1516
    wire [63:0] lut_1516_table = 64'b0000000010101010000000001010101010101010111111111010101011111111;
    wire [5:0] lut_1516_select = {
                             in_data[104],
                             in_data[9],
                             in_data[384],
                             in_data[735],
                             in_data[138],
                             in_data[636]};
    
    wire lut_1516_out = lut_1516_table[lut_1516_select];
    
    generate
    if ( USE_REG ) begin : ff_1516
        reg   lut_1516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1516_ff <= lut_1516_out;
            end
        end
        
        assign out_data[1516] = lut_1516_ff;
    end
    else begin : no_ff_1516
        assign out_data[1516] = lut_1516_out;
    end
    endgenerate
    
    
    
    // LUT : 1517
    wire [63:0] lut_1517_table = 64'b1111111111111111111111111111111101010101010101010101010101010101;
    wire [5:0] lut_1517_select = {
                             in_data[329],
                             in_data[280],
                             in_data[723],
                             in_data[56],
                             in_data[546],
                             in_data[402]};
    
    wire lut_1517_out = lut_1517_table[lut_1517_select];
    
    generate
    if ( USE_REG ) begin : ff_1517
        reg   lut_1517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1517_ff <= lut_1517_out;
            end
        end
        
        assign out_data[1517] = lut_1517_ff;
    end
    else begin : no_ff_1517
        assign out_data[1517] = lut_1517_out;
    end
    endgenerate
    
    
    
    // LUT : 1518
    wire [63:0] lut_1518_table = 64'b1111111111111111110111110101111101010101000000000100000000000000;
    wire [5:0] lut_1518_select = {
                             in_data[262],
                             in_data[535],
                             in_data[503],
                             in_data[702],
                             in_data[17],
                             in_data[445]};
    
    wire lut_1518_out = lut_1518_table[lut_1518_select];
    
    generate
    if ( USE_REG ) begin : ff_1518
        reg   lut_1518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1518_ff <= lut_1518_out;
            end
        end
        
        assign out_data[1518] = lut_1518_ff;
    end
    else begin : no_ff_1518
        assign out_data[1518] = lut_1518_out;
    end
    endgenerate
    
    
    
    // LUT : 1519
    wire [63:0] lut_1519_table = 64'b0000000000000000000000000001000000000000000000000000000011010001;
    wire [5:0] lut_1519_select = {
                             in_data[147],
                             in_data[360],
                             in_data[708],
                             in_data[638],
                             in_data[441],
                             in_data[715]};
    
    wire lut_1519_out = lut_1519_table[lut_1519_select];
    
    generate
    if ( USE_REG ) begin : ff_1519
        reg   lut_1519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1519_ff <= lut_1519_out;
            end
        end
        
        assign out_data[1519] = lut_1519_ff;
    end
    else begin : no_ff_1519
        assign out_data[1519] = lut_1519_out;
    end
    endgenerate
    
    
    
    // LUT : 1520
    wire [63:0] lut_1520_table = 64'b1111111111001111111111111100111111011111110011011101111111001101;
    wire [5:0] lut_1520_select = {
                             in_data[583],
                             in_data[141],
                             in_data[720],
                             in_data[658],
                             in_data[741],
                             in_data[70]};
    
    wire lut_1520_out = lut_1520_table[lut_1520_select];
    
    generate
    if ( USE_REG ) begin : ff_1520
        reg   lut_1520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1520_ff <= lut_1520_out;
            end
        end
        
        assign out_data[1520] = lut_1520_ff;
    end
    else begin : no_ff_1520
        assign out_data[1520] = lut_1520_out;
    end
    endgenerate
    
    
    
    // LUT : 1521
    wire [63:0] lut_1521_table = 64'b0011001100110011111111110111011100010001000000000011001100100010;
    wire [5:0] lut_1521_select = {
                             in_data[98],
                             in_data[655],
                             in_data[547],
                             in_data[335],
                             in_data[246],
                             in_data[566]};
    
    wire lut_1521_out = lut_1521_table[lut_1521_select];
    
    generate
    if ( USE_REG ) begin : ff_1521
        reg   lut_1521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1521_ff <= lut_1521_out;
            end
        end
        
        assign out_data[1521] = lut_1521_ff;
    end
    else begin : no_ff_1521
        assign out_data[1521] = lut_1521_out;
    end
    endgenerate
    
    
    
    // LUT : 1522
    wire [63:0] lut_1522_table = 64'b0000000101000000000101010100000000000001010000000000010101000000;
    wire [5:0] lut_1522_select = {
                             in_data[739],
                             in_data[746],
                             in_data[497],
                             in_data[285],
                             in_data[181],
                             in_data[690]};
    
    wire lut_1522_out = lut_1522_table[lut_1522_select];
    
    generate
    if ( USE_REG ) begin : ff_1522
        reg   lut_1522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1522_ff <= lut_1522_out;
            end
        end
        
        assign out_data[1522] = lut_1522_ff;
    end
    else begin : no_ff_1522
        assign out_data[1522] = lut_1522_out;
    end
    endgenerate
    
    
    
    // LUT : 1523
    wire [63:0] lut_1523_table = 64'b1111111111111111111111111111111110001111000011111000111010001010;
    wire [5:0] lut_1523_select = {
                             in_data[405],
                             in_data[713],
                             in_data[391],
                             in_data[630],
                             in_data[3],
                             in_data[647]};
    
    wire lut_1523_out = lut_1523_table[lut_1523_select];
    
    generate
    if ( USE_REG ) begin : ff_1523
        reg   lut_1523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1523_ff <= lut_1523_out;
            end
        end
        
        assign out_data[1523] = lut_1523_ff;
    end
    else begin : no_ff_1523
        assign out_data[1523] = lut_1523_out;
    end
    endgenerate
    
    
    
    // LUT : 1524
    wire [63:0] lut_1524_table = 64'b1011101110111011101110111011101100110011101110110011001100100010;
    wire [5:0] lut_1524_select = {
                             in_data[459],
                             in_data[595],
                             in_data[508],
                             in_data[533],
                             in_data[707],
                             in_data[686]};
    
    wire lut_1524_out = lut_1524_table[lut_1524_select];
    
    generate
    if ( USE_REG ) begin : ff_1524
        reg   lut_1524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1524_ff <= lut_1524_out;
            end
        end
        
        assign out_data[1524] = lut_1524_ff;
    end
    else begin : no_ff_1524
        assign out_data[1524] = lut_1524_out;
    end
    endgenerate
    
    
    
    // LUT : 1525
    wire [63:0] lut_1525_table = 64'b0000000000000100000000000100010000000000010001000000000001000100;
    wire [5:0] lut_1525_select = {
                             in_data[146],
                             in_data[144],
                             in_data[651],
                             in_data[757],
                             in_data[521],
                             in_data[67]};
    
    wire lut_1525_out = lut_1525_table[lut_1525_select];
    
    generate
    if ( USE_REG ) begin : ff_1525
        reg   lut_1525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1525_ff <= lut_1525_out;
            end
        end
        
        assign out_data[1525] = lut_1525_ff;
    end
    else begin : no_ff_1525
        assign out_data[1525] = lut_1525_out;
    end
    endgenerate
    
    
    
    // LUT : 1526
    wire [63:0] lut_1526_table = 64'b1110111100001100111111110000110011001111000011001111111100001100;
    wire [5:0] lut_1526_select = {
                             in_data[171],
                             in_data[47],
                             in_data[298],
                             in_data[136],
                             in_data[625],
                             in_data[38]};
    
    wire lut_1526_out = lut_1526_table[lut_1526_select];
    
    generate
    if ( USE_REG ) begin : ff_1526
        reg   lut_1526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1526_ff <= lut_1526_out;
            end
        end
        
        assign out_data[1526] = lut_1526_ff;
    end
    else begin : no_ff_1526
        assign out_data[1526] = lut_1526_out;
    end
    endgenerate
    
    
    
    // LUT : 1527
    wire [63:0] lut_1527_table = 64'b1010100010100000111110011011100110100000101100001011100110111001;
    wire [5:0] lut_1527_select = {
                             in_data[531],
                             in_data[193],
                             in_data[170],
                             in_data[303],
                             in_data[342],
                             in_data[510]};
    
    wire lut_1527_out = lut_1527_table[lut_1527_select];
    
    generate
    if ( USE_REG ) begin : ff_1527
        reg   lut_1527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1527_ff <= lut_1527_out;
            end
        end
        
        assign out_data[1527] = lut_1527_ff;
    end
    else begin : no_ff_1527
        assign out_data[1527] = lut_1527_out;
    end
    endgenerate
    
    
    
    // LUT : 1528
    wire [63:0] lut_1528_table = 64'b0010001000101010000000000000001010111011101110110010001000100010;
    wire [5:0] lut_1528_select = {
                             in_data[444],
                             in_data[202],
                             in_data[727],
                             in_data[43],
                             in_data[157],
                             in_data[490]};
    
    wire lut_1528_out = lut_1528_table[lut_1528_select];
    
    generate
    if ( USE_REG ) begin : ff_1528
        reg   lut_1528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1528_ff <= lut_1528_out;
            end
        end
        
        assign out_data[1528] = lut_1528_ff;
    end
    else begin : no_ff_1528
        assign out_data[1528] = lut_1528_out;
    end
    endgenerate
    
    
    
    // LUT : 1529
    wire [63:0] lut_1529_table = 64'b1111111111111110111111110000000011111111111010101111111100000000;
    wire [5:0] lut_1529_select = {
                             in_data[278],
                             in_data[573],
                             in_data[455],
                             in_data[694],
                             in_data[305],
                             in_data[774]};
    
    wire lut_1529_out = lut_1529_table[lut_1529_select];
    
    generate
    if ( USE_REG ) begin : ff_1529
        reg   lut_1529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1529_ff <= lut_1529_out;
            end
        end
        
        assign out_data[1529] = lut_1529_ff;
    end
    else begin : no_ff_1529
        assign out_data[1529] = lut_1529_out;
    end
    endgenerate
    
    
    
    // LUT : 1530
    wire [63:0] lut_1530_table = 64'b0000110011001100000011001100110000000100110011000000010011001100;
    wire [5:0] lut_1530_select = {
                             in_data[751],
                             in_data[142],
                             in_data[95],
                             in_data[414],
                             in_data[351],
                             in_data[542]};
    
    wire lut_1530_out = lut_1530_table[lut_1530_select];
    
    generate
    if ( USE_REG ) begin : ff_1530
        reg   lut_1530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1530_ff <= lut_1530_out;
            end
        end
        
        assign out_data[1530] = lut_1530_ff;
    end
    else begin : no_ff_1530
        assign out_data[1530] = lut_1530_out;
    end
    endgenerate
    
    
    
    // LUT : 1531
    wire [63:0] lut_1531_table = 64'b0000000000000000111100001111101000000000000000001111000011111011;
    wire [5:0] lut_1531_select = {
                             in_data[87],
                             in_data[569],
                             in_data[255],
                             in_data[234],
                             in_data[562],
                             in_data[15]};
    
    wire lut_1531_out = lut_1531_table[lut_1531_select];
    
    generate
    if ( USE_REG ) begin : ff_1531
        reg   lut_1531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1531_ff <= lut_1531_out;
            end
        end
        
        assign out_data[1531] = lut_1531_ff;
    end
    else begin : no_ff_1531
        assign out_data[1531] = lut_1531_out;
    end
    endgenerate
    
    
    
    // LUT : 1532
    wire [63:0] lut_1532_table = 64'b0000000011110101000000001111010100000000111101010000000011110101;
    wire [5:0] lut_1532_select = {
                             in_data[760],
                             in_data[502],
                             in_data[205],
                             in_data[361],
                             in_data[534],
                             in_data[327]};
    
    wire lut_1532_out = lut_1532_table[lut_1532_select];
    
    generate
    if ( USE_REG ) begin : ff_1532
        reg   lut_1532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1532_ff <= lut_1532_out;
            end
        end
        
        assign out_data[1532] = lut_1532_ff;
    end
    else begin : no_ff_1532
        assign out_data[1532] = lut_1532_out;
    end
    endgenerate
    
    
    
    // LUT : 1533
    wire [63:0] lut_1533_table = 64'b0000100000001100000000100010001000001100000011100011001100111011;
    wire [5:0] lut_1533_select = {
                             in_data[135],
                             in_data[289],
                             in_data[240],
                             in_data[626],
                             in_data[264],
                             in_data[621]};
    
    wire lut_1533_out = lut_1533_table[lut_1533_select];
    
    generate
    if ( USE_REG ) begin : ff_1533
        reg   lut_1533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1533_ff <= lut_1533_out;
            end
        end
        
        assign out_data[1533] = lut_1533_ff;
    end
    else begin : no_ff_1533
        assign out_data[1533] = lut_1533_out;
    end
    endgenerate
    
    
    
    // LUT : 1534
    wire [63:0] lut_1534_table = 64'b0011001100110011001100110000001100110011001100110011001100000011;
    wire [5:0] lut_1534_select = {
                             in_data[754],
                             in_data[680],
                             in_data[743],
                             in_data[10],
                             in_data[150],
                             in_data[449]};
    
    wire lut_1534_out = lut_1534_table[lut_1534_select];
    
    generate
    if ( USE_REG ) begin : ff_1534
        reg   lut_1534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1534_ff <= lut_1534_out;
            end
        end
        
        assign out_data[1534] = lut_1534_ff;
    end
    else begin : no_ff_1534
        assign out_data[1534] = lut_1534_out;
    end
    endgenerate
    
    
    
    // LUT : 1535
    wire [63:0] lut_1535_table = 64'b0000000000000000000000000000000000000000000000010000000000000000;
    wire [5:0] lut_1535_select = {
                             in_data[310],
                             in_data[251],
                             in_data[394],
                             in_data[766],
                             in_data[770],
                             in_data[107]};
    
    wire lut_1535_out = lut_1535_table[lut_1535_select];
    
    generate
    if ( USE_REG ) begin : ff_1535
        reg   lut_1535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1535_ff <= lut_1535_out;
            end
        end
        
        assign out_data[1535] = lut_1535_ff;
    end
    else begin : no_ff_1535
        assign out_data[1535] = lut_1535_out;
    end
    endgenerate
    
    
    
    // LUT : 1536
    wire [63:0] lut_1536_table = 64'b0000000011000000110000001111001100000000110000001100000011110011;
    wire [5:0] lut_1536_select = {
                             in_data[475],
                             in_data[71],
                             in_data[163],
                             in_data[188],
                             in_data[130],
                             in_data[674]};
    
    wire lut_1536_out = lut_1536_table[lut_1536_select];
    
    generate
    if ( USE_REG ) begin : ff_1536
        reg   lut_1536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1536_ff <= lut_1536_out;
            end
        end
        
        assign out_data[1536] = lut_1536_ff;
    end
    else begin : no_ff_1536
        assign out_data[1536] = lut_1536_out;
    end
    endgenerate
    
    
    
    // LUT : 1537
    wire [63:0] lut_1537_table = 64'b1111111111111111111111111111111111111111111111110000010000000000;
    wire [5:0] lut_1537_select = {
                             in_data[274],
                             in_data[304],
                             in_data[660],
                             in_data[65],
                             in_data[254],
                             in_data[45]};
    
    wire lut_1537_out = lut_1537_table[lut_1537_select];
    
    generate
    if ( USE_REG ) begin : ff_1537
        reg   lut_1537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1537_ff <= lut_1537_out;
            end
        end
        
        assign out_data[1537] = lut_1537_ff;
    end
    else begin : no_ff_1537
        assign out_data[1537] = lut_1537_out;
    end
    endgenerate
    
    
    
    // LUT : 1538
    wire [63:0] lut_1538_table = 64'b1111100111111000111111011111110011111111111011001111111111101000;
    wire [5:0] lut_1538_select = {
                             in_data[600],
                             in_data[652],
                             in_data[433],
                             in_data[579],
                             in_data[519],
                             in_data[124]};
    
    wire lut_1538_out = lut_1538_table[lut_1538_select];
    
    generate
    if ( USE_REG ) begin : ff_1538
        reg   lut_1538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1538_ff <= lut_1538_out;
            end
        end
        
        assign out_data[1538] = lut_1538_ff;
    end
    else begin : no_ff_1538
        assign out_data[1538] = lut_1538_out;
    end
    endgenerate
    
    
    
    // LUT : 1539
    wire [63:0] lut_1539_table = 64'b0101010101000000010101010000000011111111110111011101110101000100;
    wire [5:0] lut_1539_select = {
                             in_data[396],
                             in_data[290],
                             in_data[687],
                             in_data[756],
                             in_data[584],
                             in_data[357]};
    
    wire lut_1539_out = lut_1539_table[lut_1539_select];
    
    generate
    if ( USE_REG ) begin : ff_1539
        reg   lut_1539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1539_ff <= lut_1539_out;
            end
        end
        
        assign out_data[1539] = lut_1539_ff;
    end
    else begin : no_ff_1539
        assign out_data[1539] = lut_1539_out;
    end
    endgenerate
    
    
    
    // LUT : 1540
    wire [63:0] lut_1540_table = 64'b1111111101010101010101010101010111111111011101110101010101010101;
    wire [5:0] lut_1540_select = {
                             in_data[201],
                             in_data[632],
                             in_data[277],
                             in_data[761],
                             in_data[644],
                             in_data[239]};
    
    wire lut_1540_out = lut_1540_table[lut_1540_select];
    
    generate
    if ( USE_REG ) begin : ff_1540
        reg   lut_1540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1540_ff <= lut_1540_out;
            end
        end
        
        assign out_data[1540] = lut_1540_ff;
    end
    else begin : no_ff_1540
        assign out_data[1540] = lut_1540_out;
    end
    endgenerate
    
    
    
    // LUT : 1541
    wire [63:0] lut_1541_table = 64'b1010101011101110101010101111111110101010111011101010101011111111;
    wire [5:0] lut_1541_select = {
                             in_data[309],
                             in_data[745],
                             in_data[345],
                             in_data[587],
                             in_data[639],
                             in_data[286]};
    
    wire lut_1541_out = lut_1541_table[lut_1541_select];
    
    generate
    if ( USE_REG ) begin : ff_1541
        reg   lut_1541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1541_ff <= lut_1541_out;
            end
        end
        
        assign out_data[1541] = lut_1541_ff;
    end
    else begin : no_ff_1541
        assign out_data[1541] = lut_1541_out;
    end
    endgenerate
    
    
    
    // LUT : 1542
    wire [63:0] lut_1542_table = 64'b0000111100001111000011110000010100001111000011110000101000001010;
    wire [5:0] lut_1542_select = {
                             in_data[435],
                             in_data[256],
                             in_data[200],
                             in_data[219],
                             in_data[198],
                             in_data[688]};
    
    wire lut_1542_out = lut_1542_table[lut_1542_select];
    
    generate
    if ( USE_REG ) begin : ff_1542
        reg   lut_1542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1542_ff <= lut_1542_out;
            end
        end
        
        assign out_data[1542] = lut_1542_ff;
    end
    else begin : no_ff_1542
        assign out_data[1542] = lut_1542_out;
    end
    endgenerate
    
    
    
    // LUT : 1543
    wire [63:0] lut_1543_table = 64'b1111010111110000111111111111000011111111111111111111111111111111;
    wire [5:0] lut_1543_select = {
                             in_data[374],
                             in_data[89],
                             in_data[42],
                             in_data[668],
                             in_data[699],
                             in_data[753]};
    
    wire lut_1543_out = lut_1543_table[lut_1543_select];
    
    generate
    if ( USE_REG ) begin : ff_1543
        reg   lut_1543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1543_ff <= lut_1543_out;
            end
        end
        
        assign out_data[1543] = lut_1543_ff;
    end
    else begin : no_ff_1543
        assign out_data[1543] = lut_1543_out;
    end
    endgenerate
    
    
    
    // LUT : 1544
    wire [63:0] lut_1544_table = 64'b1110111011111110000000101111001011111110111101000100000011110000;
    wire [5:0] lut_1544_select = {
                             in_data[301],
                             in_data[358],
                             in_data[426],
                             in_data[543],
                             in_data[377],
                             in_data[443]};
    
    wire lut_1544_out = lut_1544_table[lut_1544_select];
    
    generate
    if ( USE_REG ) begin : ff_1544
        reg   lut_1544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1544_ff <= lut_1544_out;
            end
        end
        
        assign out_data[1544] = lut_1544_ff;
    end
    else begin : no_ff_1544
        assign out_data[1544] = lut_1544_out;
    end
    endgenerate
    
    
    
    // LUT : 1545
    wire [63:0] lut_1545_table = 64'b1111111111110001111111111111111111110000000000001111001011110000;
    wire [5:0] lut_1545_select = {
                             in_data[404],
                             in_data[640],
                             in_data[492],
                             in_data[663],
                             in_data[448],
                             in_data[29]};
    
    wire lut_1545_out = lut_1545_table[lut_1545_select];
    
    generate
    if ( USE_REG ) begin : ff_1545
        reg   lut_1545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1545_ff <= lut_1545_out;
            end
        end
        
        assign out_data[1545] = lut_1545_ff;
    end
    else begin : no_ff_1545
        assign out_data[1545] = lut_1545_out;
    end
    endgenerate
    
    
    
    // LUT : 1546
    wire [63:0] lut_1546_table = 64'b0000000000000000000000000000000001011111000100011111110100000000;
    wire [5:0] lut_1546_select = {
                             in_data[714],
                             in_data[215],
                             in_data[512],
                             in_data[412],
                             in_data[273],
                             in_data[149]};
    
    wire lut_1546_out = lut_1546_table[lut_1546_select];
    
    generate
    if ( USE_REG ) begin : ff_1546
        reg   lut_1546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1546_ff <= lut_1546_out;
            end
        end
        
        assign out_data[1546] = lut_1546_ff;
    end
    else begin : no_ff_1546
        assign out_data[1546] = lut_1546_out;
    end
    endgenerate
    
    
    
    // LUT : 1547
    wire [63:0] lut_1547_table = 64'b1000100010001000111011101110111010001000100010001110111011001110;
    wire [5:0] lut_1547_select = {
                             in_data[665],
                             in_data[162],
                             in_data[16],
                             in_data[111],
                             in_data[518],
                             in_data[259]};
    
    wire lut_1547_out = lut_1547_table[lut_1547_select];
    
    generate
    if ( USE_REG ) begin : ff_1547
        reg   lut_1547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1547_ff <= lut_1547_out;
            end
        end
        
        assign out_data[1547] = lut_1547_ff;
    end
    else begin : no_ff_1547
        assign out_data[1547] = lut_1547_out;
    end
    endgenerate
    
    
    
    // LUT : 1548
    wire [63:0] lut_1548_table = 64'b1111110111111101111111011111110111010101110101011101010111010101;
    wire [5:0] lut_1548_select = {
                             in_data[49],
                             in_data[223],
                             in_data[51],
                             in_data[679],
                             in_data[676],
                             in_data[370]};
    
    wire lut_1548_out = lut_1548_table[lut_1548_select];
    
    generate
    if ( USE_REG ) begin : ff_1548
        reg   lut_1548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1548_ff <= lut_1548_out;
            end
        end
        
        assign out_data[1548] = lut_1548_ff;
    end
    else begin : no_ff_1548
        assign out_data[1548] = lut_1548_out;
    end
    endgenerate
    
    
    
    // LUT : 1549
    wire [63:0] lut_1549_table = 64'b0000000000000100000000000000010000001100111111010000010011111101;
    wire [5:0] lut_1549_select = {
                             in_data[125],
                             in_data[139],
                             in_data[69],
                             in_data[325],
                             in_data[216],
                             in_data[155]};
    
    wire lut_1549_out = lut_1549_table[lut_1549_select];
    
    generate
    if ( USE_REG ) begin : ff_1549
        reg   lut_1549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1549_ff <= lut_1549_out;
            end
        end
        
        assign out_data[1549] = lut_1549_ff;
    end
    else begin : no_ff_1549
        assign out_data[1549] = lut_1549_out;
    end
    endgenerate
    
    
    
    // LUT : 1550
    wire [63:0] lut_1550_table = 64'b1010101010101010111111111111111100000000000000001111111111111111;
    wire [5:0] lut_1550_select = {
                             in_data[173],
                             in_data[599],
                             in_data[133],
                             in_data[586],
                             in_data[366],
                             in_data[321]};
    
    wire lut_1550_out = lut_1550_table[lut_1550_select];
    
    generate
    if ( USE_REG ) begin : ff_1550
        reg   lut_1550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1550_ff <= lut_1550_out;
            end
        end
        
        assign out_data[1550] = lut_1550_ff;
    end
    else begin : no_ff_1550
        assign out_data[1550] = lut_1550_out;
    end
    endgenerate
    
    
    
    // LUT : 1551
    wire [63:0] lut_1551_table = 64'b1111111111111111000000000000000011111111111111111111111101001101;
    wire [5:0] lut_1551_select = {
                             in_data[627],
                             in_data[580],
                             in_data[96],
                             in_data[773],
                             in_data[530],
                             in_data[12]};
    
    wire lut_1551_out = lut_1551_table[lut_1551_select];
    
    generate
    if ( USE_REG ) begin : ff_1551
        reg   lut_1551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1551_ff <= lut_1551_out;
            end
        end
        
        assign out_data[1551] = lut_1551_ff;
    end
    else begin : no_ff_1551
        assign out_data[1551] = lut_1551_out;
    end
    endgenerate
    
    
    
    // LUT : 1552
    wire [63:0] lut_1552_table = 64'b0111011101110111011101110111011100000000000000000000000000000000;
    wire [5:0] lut_1552_select = {
                             in_data[520],
                             in_data[113],
                             in_data[172],
                             in_data[724],
                             in_data[564],
                             in_data[189]};
    
    wire lut_1552_out = lut_1552_table[lut_1552_select];
    
    generate
    if ( USE_REG ) begin : ff_1552
        reg   lut_1552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1552_ff <= lut_1552_out;
            end
        end
        
        assign out_data[1552] = lut_1552_ff;
    end
    else begin : no_ff_1552
        assign out_data[1552] = lut_1552_out;
    end
    endgenerate
    
    
    
    // LUT : 1553
    wire [63:0] lut_1553_table = 64'b0000000000000000000000000000000001000100010101010101010001010101;
    wire [5:0] lut_1553_select = {
                             in_data[677],
                             in_data[114],
                             in_data[4],
                             in_data[2],
                             in_data[618],
                             in_data[177]};
    
    wire lut_1553_out = lut_1553_table[lut_1553_select];
    
    generate
    if ( USE_REG ) begin : ff_1553
        reg   lut_1553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1553_ff <= lut_1553_out;
            end
        end
        
        assign out_data[1553] = lut_1553_ff;
    end
    else begin : no_ff_1553
        assign out_data[1553] = lut_1553_out;
    end
    endgenerate
    
    
    
    // LUT : 1554
    wire [63:0] lut_1554_table = 64'b0000110000001100000011000000110011001111110011110000111111001111;
    wire [5:0] lut_1554_select = {
                             in_data[398],
                             in_data[420],
                             in_data[317],
                             in_data[427],
                             in_data[613],
                             in_data[26]};
    
    wire lut_1554_out = lut_1554_table[lut_1554_select];
    
    generate
    if ( USE_REG ) begin : ff_1554
        reg   lut_1554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1554_ff <= lut_1554_out;
            end
        end
        
        assign out_data[1554] = lut_1554_ff;
    end
    else begin : no_ff_1554
        assign out_data[1554] = lut_1554_out;
    end
    endgenerate
    
    
    
    // LUT : 1555
    wire [63:0] lut_1555_table = 64'b1111111100110010111111110011000011111111000000001111111100000000;
    wire [5:0] lut_1555_select = {
                             in_data[108],
                             in_data[447],
                             in_data[346],
                             in_data[684],
                             in_data[464],
                             in_data[333]};
    
    wire lut_1555_out = lut_1555_table[lut_1555_select];
    
    generate
    if ( USE_REG ) begin : ff_1555
        reg   lut_1555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1555_ff <= lut_1555_out;
            end
        end
        
        assign out_data[1555] = lut_1555_ff;
    end
    else begin : no_ff_1555
        assign out_data[1555] = lut_1555_out;
    end
    endgenerate
    
    
    
    // LUT : 1556
    wire [63:0] lut_1556_table = 64'b1111111111111111111111111111111101110101111101011101010111110101;
    wire [5:0] lut_1556_select = {
                             in_data[768],
                             in_data[693],
                             in_data[589],
                             in_data[338],
                             in_data[730],
                             in_data[631]};
    
    wire lut_1556_out = lut_1556_table[lut_1556_select];
    
    generate
    if ( USE_REG ) begin : ff_1556
        reg   lut_1556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1556_ff <= lut_1556_out;
            end
        end
        
        assign out_data[1556] = lut_1556_ff;
    end
    else begin : no_ff_1556
        assign out_data[1556] = lut_1556_out;
    end
    endgenerate
    
    
    
    // LUT : 1557
    wire [63:0] lut_1557_table = 64'b0011000000110000101100010011000100110000101100001011000110110000;
    wire [5:0] lut_1557_select = {
                             in_data[196],
                             in_data[197],
                             in_data[726],
                             in_data[253],
                             in_data[110],
                             in_data[282]};
    
    wire lut_1557_out = lut_1557_table[lut_1557_select];
    
    generate
    if ( USE_REG ) begin : ff_1557
        reg   lut_1557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1557_ff <= lut_1557_out;
            end
        end
        
        assign out_data[1557] = lut_1557_ff;
    end
    else begin : no_ff_1557
        assign out_data[1557] = lut_1557_out;
    end
    endgenerate
    
    
    
    // LUT : 1558
    wire [63:0] lut_1558_table = 64'b1111111100001111111111111010111110111111000010101111111100001010;
    wire [5:0] lut_1558_select = {
                             in_data[302],
                             in_data[670],
                             in_data[664],
                             in_data[733],
                             in_data[740],
                             in_data[222]};
    
    wire lut_1558_out = lut_1558_table[lut_1558_select];
    
    generate
    if ( USE_REG ) begin : ff_1558
        reg   lut_1558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1558_ff <= lut_1558_out;
            end
        end
        
        assign out_data[1558] = lut_1558_ff;
    end
    else begin : no_ff_1558
        assign out_data[1558] = lut_1558_out;
    end
    endgenerate
    
    
    
    // LUT : 1559
    wire [63:0] lut_1559_table = 64'b1111111111111111110010001100100011111111111111111110111011101110;
    wire [5:0] lut_1559_select = {
                             in_data[748],
                             in_data[121],
                             in_data[393],
                             in_data[728],
                             in_data[94],
                             in_data[513]};
    
    wire lut_1559_out = lut_1559_table[lut_1559_select];
    
    generate
    if ( USE_REG ) begin : ff_1559
        reg   lut_1559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1559_ff <= lut_1559_out;
            end
        end
        
        assign out_data[1559] = lut_1559_ff;
    end
    else begin : no_ff_1559
        assign out_data[1559] = lut_1559_out;
    end
    endgenerate
    
    
    
    // LUT : 1560
    wire [63:0] lut_1560_table = 64'b1010101000000000101010100000000000001010000000001010111100001000;
    wire [5:0] lut_1560_select = {
                             in_data[361],
                             in_data[145],
                             in_data[458],
                             in_data[423],
                             in_data[59],
                             in_data[429]};
    
    wire lut_1560_out = lut_1560_table[lut_1560_select];
    
    generate
    if ( USE_REG ) begin : ff_1560
        reg   lut_1560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1560_ff <= lut_1560_out;
            end
        end
        
        assign out_data[1560] = lut_1560_ff;
    end
    else begin : no_ff_1560
        assign out_data[1560] = lut_1560_out;
    end
    endgenerate
    
    
    
    // LUT : 1561
    wire [63:0] lut_1561_table = 64'b0000000000010111000000001111111100000000000000000000000000000000;
    wire [5:0] lut_1561_select = {
                             in_data[483],
                             in_data[479],
                             in_data[624],
                             in_data[41],
                             in_data[306],
                             in_data[219]};
    
    wire lut_1561_out = lut_1561_table[lut_1561_select];
    
    generate
    if ( USE_REG ) begin : ff_1561
        reg   lut_1561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1561_ff <= lut_1561_out;
            end
        end
        
        assign out_data[1561] = lut_1561_ff;
    end
    else begin : no_ff_1561
        assign out_data[1561] = lut_1561_out;
    end
    endgenerate
    
    
    
    // LUT : 1562
    wire [63:0] lut_1562_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1562_select = {
                             in_data[616],
                             in_data[401],
                             in_data[311],
                             in_data[30],
                             in_data[94],
                             in_data[776]};
    
    wire lut_1562_out = lut_1562_table[lut_1562_select];
    
    generate
    if ( USE_REG ) begin : ff_1562
        reg   lut_1562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1562_ff <= lut_1562_out;
            end
        end
        
        assign out_data[1562] = lut_1562_ff;
    end
    else begin : no_ff_1562
        assign out_data[1562] = lut_1562_out;
    end
    endgenerate
    
    
    
    // LUT : 1563
    wire [63:0] lut_1563_table = 64'b0011000000110000001100000011000000110000001100000011000000110000;
    wire [5:0] lut_1563_select = {
                             in_data[782],
                             in_data[777],
                             in_data[17],
                             in_data[544],
                             in_data[369],
                             in_data[19]};
    
    wire lut_1563_out = lut_1563_table[lut_1563_select];
    
    generate
    if ( USE_REG ) begin : ff_1563
        reg   lut_1563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1563_ff <= lut_1563_out;
            end
        end
        
        assign out_data[1563] = lut_1563_ff;
    end
    else begin : no_ff_1563
        assign out_data[1563] = lut_1563_out;
    end
    endgenerate
    
    
    
    // LUT : 1564
    wire [63:0] lut_1564_table = 64'b1100111011001000111111101110100011011110111111101111111111111110;
    wire [5:0] lut_1564_select = {
                             in_data[687],
                             in_data[195],
                             in_data[186],
                             in_data[623],
                             in_data[509],
                             in_data[621]};
    
    wire lut_1564_out = lut_1564_table[lut_1564_select];
    
    generate
    if ( USE_REG ) begin : ff_1564
        reg   lut_1564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1564_ff <= lut_1564_out;
            end
        end
        
        assign out_data[1564] = lut_1564_ff;
    end
    else begin : no_ff_1564
        assign out_data[1564] = lut_1564_out;
    end
    endgenerate
    
    
    
    // LUT : 1565
    wire [63:0] lut_1565_table = 64'b0000000000110001000000000000000000110011111101110011001100110011;
    wire [5:0] lut_1565_select = {
                             in_data[573],
                             in_data[702],
                             in_data[98],
                             in_data[20],
                             in_data[292],
                             in_data[530]};
    
    wire lut_1565_out = lut_1565_table[lut_1565_select];
    
    generate
    if ( USE_REG ) begin : ff_1565
        reg   lut_1565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1565_ff <= lut_1565_out;
            end
        end
        
        assign out_data[1565] = lut_1565_ff;
    end
    else begin : no_ff_1565
        assign out_data[1565] = lut_1565_out;
    end
    endgenerate
    
    
    
    // LUT : 1566
    wire [63:0] lut_1566_table = 64'b0000000000000000000000010001010100000000000000000001000100010101;
    wire [5:0] lut_1566_select = {
                             in_data[251],
                             in_data[596],
                             in_data[2],
                             in_data[201],
                             in_data[46],
                             in_data[202]};
    
    wire lut_1566_out = lut_1566_table[lut_1566_select];
    
    generate
    if ( USE_REG ) begin : ff_1566
        reg   lut_1566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1566_ff <= lut_1566_out;
            end
        end
        
        assign out_data[1566] = lut_1566_ff;
    end
    else begin : no_ff_1566
        assign out_data[1566] = lut_1566_out;
    end
    endgenerate
    
    
    
    // LUT : 1567
    wire [63:0] lut_1567_table = 64'b1010101110101010111111111111111110101010101010101010101010101010;
    wire [5:0] lut_1567_select = {
                             in_data[631],
                             in_data[175],
                             in_data[35],
                             in_data[25],
                             in_data[734],
                             in_data[277]};
    
    wire lut_1567_out = lut_1567_table[lut_1567_select];
    
    generate
    if ( USE_REG ) begin : ff_1567
        reg   lut_1567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1567_ff <= lut_1567_out;
            end
        end
        
        assign out_data[1567] = lut_1567_ff;
    end
    else begin : no_ff_1567
        assign out_data[1567] = lut_1567_out;
    end
    endgenerate
    
    
    
    // LUT : 1568
    wire [63:0] lut_1568_table = 64'b1111111111111111101100101011001011111111111111111011001010110010;
    wire [5:0] lut_1568_select = {
                             in_data[308],
                             in_data[484],
                             in_data[115],
                             in_data[385],
                             in_data[599],
                             in_data[93]};
    
    wire lut_1568_out = lut_1568_table[lut_1568_select];
    
    generate
    if ( USE_REG ) begin : ff_1568
        reg   lut_1568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1568_ff <= lut_1568_out;
            end
        end
        
        assign out_data[1568] = lut_1568_ff;
    end
    else begin : no_ff_1568
        assign out_data[1568] = lut_1568_out;
    end
    endgenerate
    
    
    
    // LUT : 1569
    wire [63:0] lut_1569_table = 64'b1111101100000000111111110000000011111011000000001111111100000000;
    wire [5:0] lut_1569_select = {
                             in_data[706],
                             in_data[326],
                             in_data[571],
                             in_data[12],
                             in_data[333],
                             in_data[51]};
    
    wire lut_1569_out = lut_1569_table[lut_1569_select];
    
    generate
    if ( USE_REG ) begin : ff_1569
        reg   lut_1569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1569_ff <= lut_1569_out;
            end
        end
        
        assign out_data[1569] = lut_1569_ff;
    end
    else begin : no_ff_1569
        assign out_data[1569] = lut_1569_out;
    end
    endgenerate
    
    
    
    // LUT : 1570
    wire [63:0] lut_1570_table = 64'b0000001100011011000010110000101100001011000110110000101100011011;
    wire [5:0] lut_1570_select = {
                             in_data[64],
                             in_data[135],
                             in_data[262],
                             in_data[382],
                             in_data[470],
                             in_data[400]};
    
    wire lut_1570_out = lut_1570_table[lut_1570_select];
    
    generate
    if ( USE_REG ) begin : ff_1570
        reg   lut_1570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1570_ff <= lut_1570_out;
            end
        end
        
        assign out_data[1570] = lut_1570_ff;
    end
    else begin : no_ff_1570
        assign out_data[1570] = lut_1570_out;
    end
    endgenerate
    
    
    
    // LUT : 1571
    wire [63:0] lut_1571_table = 64'b0000000100000001000000110000001100000001000000010000001100000011;
    wire [5:0] lut_1571_select = {
                             in_data[3],
                             in_data[629],
                             in_data[113],
                             in_data[412],
                             in_data[744],
                             in_data[612]};
    
    wire lut_1571_out = lut_1571_table[lut_1571_select];
    
    generate
    if ( USE_REG ) begin : ff_1571
        reg   lut_1571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1571_ff <= lut_1571_out;
            end
        end
        
        assign out_data[1571] = lut_1571_ff;
    end
    else begin : no_ff_1571
        assign out_data[1571] = lut_1571_out;
    end
    endgenerate
    
    
    
    // LUT : 1572
    wire [63:0] lut_1572_table = 64'b1111110011001100111111001100110011111100110011001111110011001100;
    wire [5:0] lut_1572_select = {
                             in_data[23],
                             in_data[18],
                             in_data[241],
                             in_data[508],
                             in_data[547],
                             in_data[672]};
    
    wire lut_1572_out = lut_1572_table[lut_1572_select];
    
    generate
    if ( USE_REG ) begin : ff_1572
        reg   lut_1572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1572_ff <= lut_1572_out;
            end
        end
        
        assign out_data[1572] = lut_1572_ff;
    end
    else begin : no_ff_1572
        assign out_data[1572] = lut_1572_out;
    end
    endgenerate
    
    
    
    // LUT : 1573
    wire [63:0] lut_1573_table = 64'b0000000011001100000000001100110000000000110011000000000011001100;
    wire [5:0] lut_1573_select = {
                             in_data[763],
                             in_data[754],
                             in_data[273],
                             in_data[578],
                             in_data[323],
                             in_data[56]};
    
    wire lut_1573_out = lut_1573_table[lut_1573_select];
    
    generate
    if ( USE_REG ) begin : ff_1573
        reg   lut_1573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1573_ff <= lut_1573_out;
            end
        end
        
        assign out_data[1573] = lut_1573_ff;
    end
    else begin : no_ff_1573
        assign out_data[1573] = lut_1573_out;
    end
    endgenerate
    
    
    
    // LUT : 1574
    wire [63:0] lut_1574_table = 64'b1010001010101011001000001010101010101010101010110010001010101010;
    wire [5:0] lut_1574_select = {
                             in_data[50],
                             in_data[194],
                             in_data[496],
                             in_data[658],
                             in_data[689],
                             in_data[295]};
    
    wire lut_1574_out = lut_1574_table[lut_1574_select];
    
    generate
    if ( USE_REG ) begin : ff_1574
        reg   lut_1574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1574_ff <= lut_1574_out;
            end
        end
        
        assign out_data[1574] = lut_1574_ff;
    end
    else begin : no_ff_1574
        assign out_data[1574] = lut_1574_out;
    end
    endgenerate
    
    
    
    // LUT : 1575
    wire [63:0] lut_1575_table = 64'b1111111111111111111111111111111111111111111111111111000011110000;
    wire [5:0] lut_1575_select = {
                             in_data[594],
                             in_data[230],
                             in_data[652],
                             in_data[575],
                             in_data[420],
                             in_data[760]};
    
    wire lut_1575_out = lut_1575_table[lut_1575_select];
    
    generate
    if ( USE_REG ) begin : ff_1575
        reg   lut_1575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1575_ff <= lut_1575_out;
            end
        end
        
        assign out_data[1575] = lut_1575_ff;
    end
    else begin : no_ff_1575
        assign out_data[1575] = lut_1575_out;
    end
    endgenerate
    
    
    
    // LUT : 1576
    wire [63:0] lut_1576_table = 64'b1111101111111111111110101111111111110000111110101010101011111010;
    wire [5:0] lut_1576_select = {
                             in_data[688],
                             in_data[417],
                             in_data[711],
                             in_data[119],
                             in_data[61],
                             in_data[579]};
    
    wire lut_1576_out = lut_1576_table[lut_1576_select];
    
    generate
    if ( USE_REG ) begin : ff_1576
        reg   lut_1576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1576_ff <= lut_1576_out;
            end
        end
        
        assign out_data[1576] = lut_1576_ff;
    end
    else begin : no_ff_1576
        assign out_data[1576] = lut_1576_out;
    end
    endgenerate
    
    
    
    // LUT : 1577
    wire [63:0] lut_1577_table = 64'b0100010001010100111111111111111100000000010000000101111101011101;
    wire [5:0] lut_1577_select = {
                             in_data[375],
                             in_data[210],
                             in_data[476],
                             in_data[74],
                             in_data[108],
                             in_data[350]};
    
    wire lut_1577_out = lut_1577_table[lut_1577_select];
    
    generate
    if ( USE_REG ) begin : ff_1577
        reg   lut_1577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1577_ff <= lut_1577_out;
            end
        end
        
        assign out_data[1577] = lut_1577_ff;
    end
    else begin : no_ff_1577
        assign out_data[1577] = lut_1577_out;
    end
    endgenerate
    
    
    
    // LUT : 1578
    wire [63:0] lut_1578_table = 64'b0101010101010101111101110111011100001101000001010011000000010001;
    wire [5:0] lut_1578_select = {
                             in_data[684],
                             in_data[246],
                             in_data[71],
                             in_data[461],
                             in_data[467],
                             in_data[220]};
    
    wire lut_1578_out = lut_1578_table[lut_1578_select];
    
    generate
    if ( USE_REG ) begin : ff_1578
        reg   lut_1578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1578_ff <= lut_1578_out;
            end
        end
        
        assign out_data[1578] = lut_1578_ff;
    end
    else begin : no_ff_1578
        assign out_data[1578] = lut_1578_out;
    end
    endgenerate
    
    
    
    // LUT : 1579
    wire [63:0] lut_1579_table = 64'b1111101011111010111110101111101011111010111110101111101011111010;
    wire [5:0] lut_1579_select = {
                             in_data[162],
                             in_data[24],
                             in_data[112],
                             in_data[635],
                             in_data[114],
                             in_data[433]};
    
    wire lut_1579_out = lut_1579_table[lut_1579_select];
    
    generate
    if ( USE_REG ) begin : ff_1579
        reg   lut_1579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1579_ff <= lut_1579_out;
            end
        end
        
        assign out_data[1579] = lut_1579_ff;
    end
    else begin : no_ff_1579
        assign out_data[1579] = lut_1579_out;
    end
    endgenerate
    
    
    
    // LUT : 1580
    wire [63:0] lut_1580_table = 64'b0100010101010101000000000000000011111111111111110000000000000000;
    wire [5:0] lut_1580_select = {
                             in_data[442],
                             in_data[294],
                             in_data[44],
                             in_data[590],
                             in_data[653],
                             in_data[208]};
    
    wire lut_1580_out = lut_1580_table[lut_1580_select];
    
    generate
    if ( USE_REG ) begin : ff_1580
        reg   lut_1580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1580_ff <= lut_1580_out;
            end
        end
        
        assign out_data[1580] = lut_1580_ff;
    end
    else begin : no_ff_1580
        assign out_data[1580] = lut_1580_out;
    end
    endgenerate
    
    
    
    // LUT : 1581
    wire [63:0] lut_1581_table = 64'b0000000000001000000000000000000000001111000011110000000000001100;
    wire [5:0] lut_1581_select = {
                             in_data[667],
                             in_data[690],
                             in_data[415],
                             in_data[565],
                             in_data[318],
                             in_data[533]};
    
    wire lut_1581_out = lut_1581_table[lut_1581_select];
    
    generate
    if ( USE_REG ) begin : ff_1581
        reg   lut_1581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1581_ff <= lut_1581_out;
            end
        end
        
        assign out_data[1581] = lut_1581_ff;
    end
    else begin : no_ff_1581
        assign out_data[1581] = lut_1581_out;
    end
    endgenerate
    
    
    
    // LUT : 1582
    wire [63:0] lut_1582_table = 64'b1111000000000000111111111111111111100000000000001010000010101110;
    wire [5:0] lut_1582_select = {
                             in_data[177],
                             in_data[218],
                             in_data[324],
                             in_data[298],
                             in_data[171],
                             in_data[602]};
    
    wire lut_1582_out = lut_1582_table[lut_1582_select];
    
    generate
    if ( USE_REG ) begin : ff_1582
        reg   lut_1582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1582_ff <= lut_1582_out;
            end
        end
        
        assign out_data[1582] = lut_1582_ff;
    end
    else begin : no_ff_1582
        assign out_data[1582] = lut_1582_out;
    end
    endgenerate
    
    
    
    // LUT : 1583
    wire [63:0] lut_1583_table = 64'b1111111111111111111111111111111111111111111111111111111011111110;
    wire [5:0] lut_1583_select = {
                             in_data[284],
                             in_data[69],
                             in_data[729],
                             in_data[79],
                             in_data[172],
                             in_data[192]};
    
    wire lut_1583_out = lut_1583_table[lut_1583_select];
    
    generate
    if ( USE_REG ) begin : ff_1583
        reg   lut_1583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1583_ff <= lut_1583_out;
            end
        end
        
        assign out_data[1583] = lut_1583_ff;
    end
    else begin : no_ff_1583
        assign out_data[1583] = lut_1583_out;
    end
    endgenerate
    
    
    
    // LUT : 1584
    wire [63:0] lut_1584_table = 64'b1111111111111111111111001111110011111111111111101111110011111100;
    wire [5:0] lut_1584_select = {
                             in_data[88],
                             in_data[258],
                             in_data[719],
                             in_data[329],
                             in_data[746],
                             in_data[16]};
    
    wire lut_1584_out = lut_1584_table[lut_1584_select];
    
    generate
    if ( USE_REG ) begin : ff_1584
        reg   lut_1584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1584_ff <= lut_1584_out;
            end
        end
        
        assign out_data[1584] = lut_1584_ff;
    end
    else begin : no_ff_1584
        assign out_data[1584] = lut_1584_out;
    end
    endgenerate
    
    
    
    // LUT : 1585
    wire [63:0] lut_1585_table = 64'b0000000000000000000000000100010001000100010001000100010001010100;
    wire [5:0] lut_1585_select = {
                             in_data[693],
                             in_data[506],
                             in_data[769],
                             in_data[362],
                             in_data[510],
                             in_data[148]};
    
    wire lut_1585_out = lut_1585_table[lut_1585_select];
    
    generate
    if ( USE_REG ) begin : ff_1585
        reg   lut_1585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1585_ff <= lut_1585_out;
            end
        end
        
        assign out_data[1585] = lut_1585_ff;
    end
    else begin : no_ff_1585
        assign out_data[1585] = lut_1585_out;
    end
    endgenerate
    
    
    
    // LUT : 1586
    wire [63:0] lut_1586_table = 64'b1000100011001000111111111111111100000000010001001101110111011111;
    wire [5:0] lut_1586_select = {
                             in_data[331],
                             in_data[185],
                             in_data[110],
                             in_data[252],
                             in_data[193],
                             in_data[538]};
    
    wire lut_1586_out = lut_1586_table[lut_1586_select];
    
    generate
    if ( USE_REG ) begin : ff_1586
        reg   lut_1586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1586_ff <= lut_1586_out;
            end
        end
        
        assign out_data[1586] = lut_1586_ff;
    end
    else begin : no_ff_1586
        assign out_data[1586] = lut_1586_out;
    end
    endgenerate
    
    
    
    // LUT : 1587
    wire [63:0] lut_1587_table = 64'b0000000000100000111111111111011100000000000000001111111101110101;
    wire [5:0] lut_1587_select = {
                             in_data[222],
                             in_data[272],
                             in_data[131],
                             in_data[526],
                             in_data[450],
                             in_data[516]};
    
    wire lut_1587_out = lut_1587_table[lut_1587_select];
    
    generate
    if ( USE_REG ) begin : ff_1587
        reg   lut_1587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1587_ff <= lut_1587_out;
            end
        end
        
        assign out_data[1587] = lut_1587_ff;
    end
    else begin : no_ff_1587
        assign out_data[1587] = lut_1587_out;
    end
    endgenerate
    
    
    
    // LUT : 1588
    wire [63:0] lut_1588_table = 64'b1111000011110000000000000000000011110000111100000000000011110000;
    wire [5:0] lut_1588_select = {
                             in_data[717],
                             in_data[356],
                             in_data[680],
                             in_data[541],
                             in_data[15],
                             in_data[170]};
    
    wire lut_1588_out = lut_1588_table[lut_1588_select];
    
    generate
    if ( USE_REG ) begin : ff_1588
        reg   lut_1588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1588_ff <= lut_1588_out;
            end
        end
        
        assign out_data[1588] = lut_1588_ff;
    end
    else begin : no_ff_1588
        assign out_data[1588] = lut_1588_out;
    end
    endgenerate
    
    
    
    // LUT : 1589
    wire [63:0] lut_1589_table = 64'b0000000000100010001000100010001000000000001000100010001000100010;
    wire [5:0] lut_1589_select = {
                             in_data[728],
                             in_data[739],
                             in_data[619],
                             in_data[392],
                             in_data[99],
                             in_data[235]};
    
    wire lut_1589_out = lut_1589_table[lut_1589_select];
    
    generate
    if ( USE_REG ) begin : ff_1589
        reg   lut_1589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1589_ff <= lut_1589_out;
            end
        end
        
        assign out_data[1589] = lut_1589_ff;
    end
    else begin : no_ff_1589
        assign out_data[1589] = lut_1589_out;
    end
    endgenerate
    
    
    
    // LUT : 1590
    wire [63:0] lut_1590_table = 64'b0000000000000000000000000000000011110000011100001111011111111111;
    wire [5:0] lut_1590_select = {
                             in_data[248],
                             in_data[465],
                             in_data[39],
                             in_data[472],
                             in_data[389],
                             in_data[77]};
    
    wire lut_1590_out = lut_1590_table[lut_1590_select];
    
    generate
    if ( USE_REG ) begin : ff_1590
        reg   lut_1590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1590_ff <= lut_1590_out;
            end
        end
        
        assign out_data[1590] = lut_1590_ff;
    end
    else begin : no_ff_1590
        assign out_data[1590] = lut_1590_out;
    end
    endgenerate
    
    
    
    // LUT : 1591
    wire [63:0] lut_1591_table = 64'b1111111111111111111111111111111110101010101010100000000000000000;
    wire [5:0] lut_1591_select = {
                             in_data[268],
                             in_data[123],
                             in_data[474],
                             in_data[363],
                             in_data[699],
                             in_data[683]};
    
    wire lut_1591_out = lut_1591_table[lut_1591_select];
    
    generate
    if ( USE_REG ) begin : ff_1591
        reg   lut_1591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1591_ff <= lut_1591_out;
            end
        end
        
        assign out_data[1591] = lut_1591_ff;
    end
    else begin : no_ff_1591
        assign out_data[1591] = lut_1591_out;
    end
    endgenerate
    
    
    
    // LUT : 1592
    wire [63:0] lut_1592_table = 64'b1111111100100010111111110010001011111111001000101011111100101010;
    wire [5:0] lut_1592_select = {
                             in_data[640],
                             in_data[752],
                             in_data[95],
                             in_data[165],
                             in_data[625],
                             in_data[439]};
    
    wire lut_1592_out = lut_1592_table[lut_1592_select];
    
    generate
    if ( USE_REG ) begin : ff_1592
        reg   lut_1592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1592_ff <= lut_1592_out;
            end
        end
        
        assign out_data[1592] = lut_1592_ff;
    end
    else begin : no_ff_1592
        assign out_data[1592] = lut_1592_out;
    end
    endgenerate
    
    
    
    // LUT : 1593
    wire [63:0] lut_1593_table = 64'b0000000010111011000000101011111100000000101110110000001010111111;
    wire [5:0] lut_1593_select = {
                             in_data[477],
                             in_data[471],
                             in_data[462],
                             in_data[444],
                             in_data[68],
                             in_data[593]};
    
    wire lut_1593_out = lut_1593_table[lut_1593_select];
    
    generate
    if ( USE_REG ) begin : ff_1593
        reg   lut_1593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1593_ff <= lut_1593_out;
            end
        end
        
        assign out_data[1593] = lut_1593_ff;
    end
    else begin : no_ff_1593
        assign out_data[1593] = lut_1593_out;
    end
    endgenerate
    
    
    
    // LUT : 1594
    wire [63:0] lut_1594_table = 64'b1111111000100000101010000000000011111111101111111111111100100000;
    wire [5:0] lut_1594_select = {
                             in_data[708],
                             in_data[75],
                             in_data[490],
                             in_data[542],
                             in_data[128],
                             in_data[430]};
    
    wire lut_1594_out = lut_1594_table[lut_1594_select];
    
    generate
    if ( USE_REG ) begin : ff_1594
        reg   lut_1594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1594_ff <= lut_1594_out;
            end
        end
        
        assign out_data[1594] = lut_1594_ff;
    end
    else begin : no_ff_1594
        assign out_data[1594] = lut_1594_out;
    end
    endgenerate
    
    
    
    // LUT : 1595
    wire [63:0] lut_1595_table = 64'b1111111111111111000000001010001000000000111111110000000000000000;
    wire [5:0] lut_1595_select = {
                             in_data[481],
                             in_data[428],
                             in_data[722],
                             in_data[48],
                             in_data[419],
                             in_data[505]};
    
    wire lut_1595_out = lut_1595_table[lut_1595_select];
    
    generate
    if ( USE_REG ) begin : ff_1595
        reg   lut_1595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1595_ff <= lut_1595_out;
            end
        end
        
        assign out_data[1595] = lut_1595_ff;
    end
    else begin : no_ff_1595
        assign out_data[1595] = lut_1595_out;
    end
    endgenerate
    
    
    
    // LUT : 1596
    wire [63:0] lut_1596_table = 64'b1111111111001111111111111111111111001100110011001100000011000000;
    wire [5:0] lut_1596_select = {
                             in_data[156],
                             in_data[213],
                             in_data[552],
                             in_data[545],
                             in_data[554],
                             in_data[223]};
    
    wire lut_1596_out = lut_1596_table[lut_1596_select];
    
    generate
    if ( USE_REG ) begin : ff_1596
        reg   lut_1596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1596_ff <= lut_1596_out;
            end
        end
        
        assign out_data[1596] = lut_1596_ff;
    end
    else begin : no_ff_1596
        assign out_data[1596] = lut_1596_out;
    end
    endgenerate
    
    
    
    // LUT : 1597
    wire [63:0] lut_1597_table = 64'b1111111111111111111110101111101011111111111111111111001011111011;
    wire [5:0] lut_1597_select = {
                             in_data[205],
                             in_data[397],
                             in_data[559],
                             in_data[709],
                             in_data[287],
                             in_data[257]};
    
    wire lut_1597_out = lut_1597_table[lut_1597_select];
    
    generate
    if ( USE_REG ) begin : ff_1597
        reg   lut_1597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1597_ff <= lut_1597_out;
            end
        end
        
        assign out_data[1597] = lut_1597_ff;
    end
    else begin : no_ff_1597
        assign out_data[1597] = lut_1597_out;
    end
    endgenerate
    
    
    
    // LUT : 1598
    wire [63:0] lut_1598_table = 64'b0000101000001010111111111111111100001000000010101111111111111111;
    wire [5:0] lut_1598_select = {
                             in_data[58],
                             in_data[574],
                             in_data[336],
                             in_data[637],
                             in_data[727],
                             in_data[190]};
    
    wire lut_1598_out = lut_1598_table[lut_1598_select];
    
    generate
    if ( USE_REG ) begin : ff_1598
        reg   lut_1598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1598_ff <= lut_1598_out;
            end
        end
        
        assign out_data[1598] = lut_1598_ff;
    end
    else begin : no_ff_1598
        assign out_data[1598] = lut_1598_out;
    end
    endgenerate
    
    
    
    // LUT : 1599
    wire [63:0] lut_1599_table = 64'b1111010001000100111111011111110111110100110001001111110111111101;
    wire [5:0] lut_1599_select = {
                             in_data[55],
                             in_data[633],
                             in_data[601],
                             in_data[314],
                             in_data[564],
                             in_data[632]};
    
    wire lut_1599_out = lut_1599_table[lut_1599_select];
    
    generate
    if ( USE_REG ) begin : ff_1599
        reg   lut_1599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1599_ff <= lut_1599_out;
            end
        end
        
        assign out_data[1599] = lut_1599_ff;
    end
    else begin : no_ff_1599
        assign out_data[1599] = lut_1599_out;
    end
    endgenerate
    
    
    
    // LUT : 1600
    wire [63:0] lut_1600_table = 64'b1111011111111111111111111111111100000000000000000000000010111111;
    wire [5:0] lut_1600_select = {
                             in_data[676],
                             in_data[749],
                             in_data[704],
                             in_data[9],
                             in_data[0],
                             in_data[503]};
    
    wire lut_1600_out = lut_1600_table[lut_1600_select];
    
    generate
    if ( USE_REG ) begin : ff_1600
        reg   lut_1600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1600_ff <= lut_1600_out;
            end
        end
        
        assign out_data[1600] = lut_1600_ff;
    end
    else begin : no_ff_1600
        assign out_data[1600] = lut_1600_out;
    end
    endgenerate
    
    
    
    // LUT : 1601
    wire [63:0] lut_1601_table = 64'b0000000000001111000011001100111100000000000011000000000000001100;
    wire [5:0] lut_1601_select = {
                             in_data[182],
                             in_data[76],
                             in_data[585],
                             in_data[620],
                             in_data[231],
                             in_data[34]};
    
    wire lut_1601_out = lut_1601_table[lut_1601_select];
    
    generate
    if ( USE_REG ) begin : ff_1601
        reg   lut_1601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1601_ff <= lut_1601_out;
            end
        end
        
        assign out_data[1601] = lut_1601_ff;
    end
    else begin : no_ff_1601
        assign out_data[1601] = lut_1601_out;
    end
    endgenerate
    
    
    
    // LUT : 1602
    wire [63:0] lut_1602_table = 64'b0000000000010101000000110011111100000000000000000001000000010101;
    wire [5:0] lut_1602_select = {
                             in_data[469],
                             in_data[611],
                             in_data[413],
                             in_data[453],
                             in_data[372],
                             in_data[740]};
    
    wire lut_1602_out = lut_1602_table[lut_1602_select];
    
    generate
    if ( USE_REG ) begin : ff_1602
        reg   lut_1602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1602_ff <= lut_1602_out;
            end
        end
        
        assign out_data[1602] = lut_1602_ff;
    end
    else begin : no_ff_1602
        assign out_data[1602] = lut_1602_out;
    end
    endgenerate
    
    
    
    // LUT : 1603
    wire [63:0] lut_1603_table = 64'b1111111111111111111111111111111111111110111011101010101010101010;
    wire [5:0] lut_1603_select = {
                             in_data[340],
                             in_data[214],
                             in_data[26],
                             in_data[644],
                             in_data[626],
                             in_data[288]};
    
    wire lut_1603_out = lut_1603_table[lut_1603_select];
    
    generate
    if ( USE_REG ) begin : ff_1603
        reg   lut_1603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1603_ff <= lut_1603_out;
            end
        end
        
        assign out_data[1603] = lut_1603_ff;
    end
    else begin : no_ff_1603
        assign out_data[1603] = lut_1603_out;
    end
    endgenerate
    
    
    
    // LUT : 1604
    wire [63:0] lut_1604_table = 64'b0000000000000000110011101110111100000000000010001100111011101111;
    wire [5:0] lut_1604_select = {
                             in_data[167],
                             in_data[358],
                             in_data[399],
                             in_data[759],
                             in_data[151],
                             in_data[116]};
    
    wire lut_1604_out = lut_1604_table[lut_1604_select];
    
    generate
    if ( USE_REG ) begin : ff_1604
        reg   lut_1604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1604_ff <= lut_1604_out;
            end
        end
        
        assign out_data[1604] = lut_1604_ff;
    end
    else begin : no_ff_1604
        assign out_data[1604] = lut_1604_out;
    end
    endgenerate
    
    
    
    // LUT : 1605
    wire [63:0] lut_1605_table = 64'b1101110111111111110111011111111100000000111010100000000010001000;
    wire [5:0] lut_1605_select = {
                             in_data[431],
                             in_data[485],
                             in_data[325],
                             in_data[446],
                             in_data[405],
                             in_data[158]};
    
    wire lut_1605_out = lut_1605_table[lut_1605_select];
    
    generate
    if ( USE_REG ) begin : ff_1605
        reg   lut_1605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1605_ff <= lut_1605_out;
            end
        end
        
        assign out_data[1605] = lut_1605_ff;
    end
    else begin : no_ff_1605
        assign out_data[1605] = lut_1605_out;
    end
    endgenerate
    
    
    
    // LUT : 1606
    wire [63:0] lut_1606_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_1606_select = {
                             in_data[528],
                             in_data[313],
                             in_data[216],
                             in_data[54],
                             in_data[562],
                             in_data[337]};
    
    wire lut_1606_out = lut_1606_table[lut_1606_select];
    
    generate
    if ( USE_REG ) begin : ff_1606
        reg   lut_1606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1606_ff <= lut_1606_out;
            end
        end
        
        assign out_data[1606] = lut_1606_ff;
    end
    else begin : no_ff_1606
        assign out_data[1606] = lut_1606_out;
    end
    endgenerate
    
    
    
    // LUT : 1607
    wire [63:0] lut_1607_table = 64'b0000000000000000110111011111111100000000000000000101000101010111;
    wire [5:0] lut_1607_select = {
                             in_data[714],
                             in_data[343],
                             in_data[357],
                             in_data[37],
                             in_data[495],
                             in_data[259]};
    
    wire lut_1607_out = lut_1607_table[lut_1607_select];
    
    generate
    if ( USE_REG ) begin : ff_1607
        reg   lut_1607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1607_ff <= lut_1607_out;
            end
        end
        
        assign out_data[1607] = lut_1607_ff;
    end
    else begin : no_ff_1607
        assign out_data[1607] = lut_1607_out;
    end
    endgenerate
    
    
    
    // LUT : 1608
    wire [63:0] lut_1608_table = 64'b1111000011110000111100001111000011111011111110111111000111111001;
    wire [5:0] lut_1608_select = {
                             in_data[179],
                             in_data[364],
                             in_data[502],
                             in_data[341],
                             in_data[66],
                             in_data[398]};
    
    wire lut_1608_out = lut_1608_table[lut_1608_select];
    
    generate
    if ( USE_REG ) begin : ff_1608
        reg   lut_1608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1608_ff <= lut_1608_out;
            end
        end
        
        assign out_data[1608] = lut_1608_ff;
    end
    else begin : no_ff_1608
        assign out_data[1608] = lut_1608_out;
    end
    endgenerate
    
    
    
    // LUT : 1609
    wire [63:0] lut_1609_table = 64'b1111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_1609_select = {
                             in_data[383],
                             in_data[111],
                             in_data[240],
                             in_data[316],
                             in_data[768],
                             in_data[523]};
    
    wire lut_1609_out = lut_1609_table[lut_1609_select];
    
    generate
    if ( USE_REG ) begin : ff_1609
        reg   lut_1609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1609_ff <= lut_1609_out;
            end
        end
        
        assign out_data[1609] = lut_1609_ff;
    end
    else begin : no_ff_1609
        assign out_data[1609] = lut_1609_out;
    end
    endgenerate
    
    
    
    // LUT : 1610
    wire [63:0] lut_1610_table = 64'b0000000000000000000100010001000100000000000000000001000100010001;
    wire [5:0] lut_1610_select = {
                             in_data[677],
                             in_data[608],
                             in_data[780],
                             in_data[166],
                             in_data[126],
                             in_data[525]};
    
    wire lut_1610_out = lut_1610_table[lut_1610_select];
    
    generate
    if ( USE_REG ) begin : ff_1610
        reg   lut_1610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1610_ff <= lut_1610_out;
            end
        end
        
        assign out_data[1610] = lut_1610_ff;
    end
    else begin : no_ff_1610
        assign out_data[1610] = lut_1610_out;
    end
    endgenerate
    
    
    
    // LUT : 1611
    wire [63:0] lut_1611_table = 64'b0011001100100011001100110010001100110011001000110011001100000011;
    wire [5:0] lut_1611_select = {
                             in_data[281],
                             in_data[141],
                             in_data[432],
                             in_data[500],
                             in_data[551],
                             in_data[697]};
    
    wire lut_1611_out = lut_1611_table[lut_1611_select];
    
    generate
    if ( USE_REG ) begin : ff_1611
        reg   lut_1611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1611_ff <= lut_1611_out;
            end
        end
        
        assign out_data[1611] = lut_1611_ff;
    end
    else begin : no_ff_1611
        assign out_data[1611] = lut_1611_out;
    end
    endgenerate
    
    
    
    // LUT : 1612
    wire [63:0] lut_1612_table = 64'b0000000000000000000000000000000010111011111111111010101011111111;
    wire [5:0] lut_1612_select = {
                             in_data[406],
                             in_data[52],
                             in_data[441],
                             in_data[212],
                             in_data[418],
                             in_data[342]};
    
    wire lut_1612_out = lut_1612_table[lut_1612_select];
    
    generate
    if ( USE_REG ) begin : ff_1612
        reg   lut_1612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1612_ff <= lut_1612_out;
            end
        end
        
        assign out_data[1612] = lut_1612_ff;
    end
    else begin : no_ff_1612
        assign out_data[1612] = lut_1612_out;
    end
    endgenerate
    
    
    
    // LUT : 1613
    wire [63:0] lut_1613_table = 64'b0100010101000101000101110001011111001100110011000100110001001100;
    wire [5:0] lut_1613_select = {
                             in_data[402],
                             in_data[243],
                             in_data[733],
                             in_data[660],
                             in_data[376],
                             in_data[249]};
    
    wire lut_1613_out = lut_1613_table[lut_1613_select];
    
    generate
    if ( USE_REG ) begin : ff_1613
        reg   lut_1613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1613_ff <= lut_1613_out;
            end
        end
        
        assign out_data[1613] = lut_1613_ff;
    end
    else begin : no_ff_1613
        assign out_data[1613] = lut_1613_out;
    end
    endgenerate
    
    
    
    // LUT : 1614
    wire [63:0] lut_1614_table = 64'b0000000001010000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_1614_select = {
                             in_data[373],
                             in_data[591],
                             in_data[206],
                             in_data[524],
                             in_data[449],
                             in_data[577]};
    
    wire lut_1614_out = lut_1614_table[lut_1614_select];
    
    generate
    if ( USE_REG ) begin : ff_1614
        reg   lut_1614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1614_ff <= lut_1614_out;
            end
        end
        
        assign out_data[1614] = lut_1614_ff;
    end
    else begin : no_ff_1614
        assign out_data[1614] = lut_1614_out;
    end
    endgenerate
    
    
    
    // LUT : 1615
    wire [63:0] lut_1615_table = 64'b1100110011001100110011001100110011111100111111011110110011111101;
    wire [5:0] lut_1615_select = {
                             in_data[741],
                             in_data[671],
                             in_data[327],
                             in_data[106],
                             in_data[582],
                             in_data[774]};
    
    wire lut_1615_out = lut_1615_table[lut_1615_select];
    
    generate
    if ( USE_REG ) begin : ff_1615
        reg   lut_1615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1615_ff <= lut_1615_out;
            end
        end
        
        assign out_data[1615] = lut_1615_ff;
    end
    else begin : no_ff_1615
        assign out_data[1615] = lut_1615_out;
    end
    endgenerate
    
    
    
    // LUT : 1616
    wire [63:0] lut_1616_table = 64'b0000000000000000111111111111111111111111000000001111111101011111;
    wire [5:0] lut_1616_select = {
                             in_data[600],
                             in_data[297],
                             in_data[691],
                             in_data[642],
                             in_data[448],
                             in_data[32]};
    
    wire lut_1616_out = lut_1616_table[lut_1616_select];
    
    generate
    if ( USE_REG ) begin : ff_1616
        reg   lut_1616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1616_ff <= lut_1616_out;
            end
        end
        
        assign out_data[1616] = lut_1616_ff;
    end
    else begin : no_ff_1616
        assign out_data[1616] = lut_1616_out;
    end
    endgenerate
    
    
    
    // LUT : 1617
    wire [63:0] lut_1617_table = 64'b1101010111010101110101011101110111011101110111011101010111011101;
    wire [5:0] lut_1617_select = {
                             in_data[557],
                             in_data[90],
                             in_data[63],
                             in_data[685],
                             in_data[207],
                             in_data[520]};
    
    wire lut_1617_out = lut_1617_table[lut_1617_select];
    
    generate
    if ( USE_REG ) begin : ff_1617
        reg   lut_1617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1617_ff <= lut_1617_out;
            end
        end
        
        assign out_data[1617] = lut_1617_ff;
    end
    else begin : no_ff_1617
        assign out_data[1617] = lut_1617_out;
    end
    endgenerate
    
    
    
    // LUT : 1618
    wire [63:0] lut_1618_table = 64'b0000110000000000000000001111010000000000000000000000000011111111;
    wire [5:0] lut_1618_select = {
                             in_data[519],
                             in_data[657],
                             in_data[659],
                             in_data[348],
                             in_data[28],
                             in_data[773]};
    
    wire lut_1618_out = lut_1618_table[lut_1618_select];
    
    generate
    if ( USE_REG ) begin : ff_1618
        reg   lut_1618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1618_ff <= lut_1618_out;
            end
        end
        
        assign out_data[1618] = lut_1618_ff;
    end
    else begin : no_ff_1618
        assign out_data[1618] = lut_1618_out;
    end
    endgenerate
    
    
    
    // LUT : 1619
    wire [63:0] lut_1619_table = 64'b1011101110111011101010101010101010111010101110100010101000101010;
    wire [5:0] lut_1619_select = {
                             in_data[330],
                             in_data[265],
                             in_data[280],
                             in_data[558],
                             in_data[404],
                             in_data[346]};
    
    wire lut_1619_out = lut_1619_table[lut_1619_select];
    
    generate
    if ( USE_REG ) begin : ff_1619
        reg   lut_1619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1619_ff <= lut_1619_out;
            end
        end
        
        assign out_data[1619] = lut_1619_ff;
    end
    else begin : no_ff_1619
        assign out_data[1619] = lut_1619_out;
    end
    endgenerate
    
    
    
    // LUT : 1620
    wire [63:0] lut_1620_table = 64'b0101010101010101010101011111110101010000111101010101000011110101;
    wire [5:0] lut_1620_select = {
                             in_data[187],
                             in_data[322],
                             in_data[745],
                             in_data[315],
                             in_data[767],
                             in_data[238]};
    
    wire lut_1620_out = lut_1620_table[lut_1620_select];
    
    generate
    if ( USE_REG ) begin : ff_1620
        reg   lut_1620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1620_ff <= lut_1620_out;
            end
        end
        
        assign out_data[1620] = lut_1620_ff;
    end
    else begin : no_ff_1620
        assign out_data[1620] = lut_1620_out;
    end
    endgenerate
    
    
    
    // LUT : 1621
    wire [63:0] lut_1621_table = 64'b1000100000000000110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1621_select = {
                             in_data[713],
                             in_data[724],
                             in_data[645],
                             in_data[45],
                             in_data[411],
                             in_data[225]};
    
    wire lut_1621_out = lut_1621_table[lut_1621_select];
    
    generate
    if ( USE_REG ) begin : ff_1621
        reg   lut_1621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1621_ff <= lut_1621_out;
            end
        end
        
        assign out_data[1621] = lut_1621_ff;
    end
    else begin : no_ff_1621
        assign out_data[1621] = lut_1621_out;
    end
    endgenerate
    
    
    
    // LUT : 1622
    wire [63:0] lut_1622_table = 64'b0000111000001101111111111101110100001110000000001110111100001100;
    wire [5:0] lut_1622_select = {
                             in_data[275],
                             in_data[598],
                             in_data[517],
                             in_data[679],
                             in_data[636],
                             in_data[233]};
    
    wire lut_1622_out = lut_1622_table[lut_1622_select];
    
    generate
    if ( USE_REG ) begin : ff_1622
        reg   lut_1622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1622_ff <= lut_1622_out;
            end
        end
        
        assign out_data[1622] = lut_1622_ff;
    end
    else begin : no_ff_1622
        assign out_data[1622] = lut_1622_out;
    end
    endgenerate
    
    
    
    // LUT : 1623
    wire [63:0] lut_1623_table = 64'b0000000000000000000000000000000000000000111111110000000011111111;
    wire [5:0] lut_1623_select = {
                             in_data[217],
                             in_data[228],
                             in_data[101],
                             in_data[390],
                             in_data[549],
                             in_data[84]};
    
    wire lut_1623_out = lut_1623_table[lut_1623_select];
    
    generate
    if ( USE_REG ) begin : ff_1623
        reg   lut_1623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1623_ff <= lut_1623_out;
            end
        end
        
        assign out_data[1623] = lut_1623_ff;
    end
    else begin : no_ff_1623
        assign out_data[1623] = lut_1623_out;
    end
    endgenerate
    
    
    
    // LUT : 1624
    wire [63:0] lut_1624_table = 64'b0000000000000000000000000000000000000000000000110000001100000011;
    wire [5:0] lut_1624_select = {
                             in_data[497],
                             in_data[253],
                             in_data[1],
                             in_data[537],
                             in_data[414],
                             in_data[60]};
    
    wire lut_1624_out = lut_1624_table[lut_1624_select];
    
    generate
    if ( USE_REG ) begin : ff_1624
        reg   lut_1624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1624_ff <= lut_1624_out;
            end
        end
        
        assign out_data[1624] = lut_1624_ff;
    end
    else begin : no_ff_1624
        assign out_data[1624] = lut_1624_out;
    end
    endgenerate
    
    
    
    // LUT : 1625
    wire [63:0] lut_1625_table = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    wire [5:0] lut_1625_select = {
                             in_data[675],
                             in_data[105],
                             in_data[319],
                             in_data[200],
                             in_data[255],
                             in_data[589]};
    
    wire lut_1625_out = lut_1625_table[lut_1625_select];
    
    generate
    if ( USE_REG ) begin : ff_1625
        reg   lut_1625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1625_ff <= lut_1625_out;
            end
        end
        
        assign out_data[1625] = lut_1625_ff;
    end
    else begin : no_ff_1625
        assign out_data[1625] = lut_1625_out;
    end
    endgenerate
    
    
    
    // LUT : 1626
    wire [63:0] lut_1626_table = 64'b1111111100000101111110110000000000001010000001011111111100000101;
    wire [5:0] lut_1626_select = {
                             in_data[664],
                             in_data[153],
                             in_data[597],
                             in_data[661],
                             in_data[617],
                             in_data[134]};
    
    wire lut_1626_out = lut_1626_table[lut_1626_select];
    
    generate
    if ( USE_REG ) begin : ff_1626
        reg   lut_1626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1626_ff <= lut_1626_out;
            end
        end
        
        assign out_data[1626] = lut_1626_ff;
    end
    else begin : no_ff_1626
        assign out_data[1626] = lut_1626_out;
    end
    endgenerate
    
    
    
    // LUT : 1627
    wire [63:0] lut_1627_table = 64'b0101010100000100010101010000010001010101000000000101010100000000;
    wire [5:0] lut_1627_select = {
                             in_data[535],
                             in_data[532],
                             in_data[211],
                             in_data[197],
                             in_data[723],
                             in_data[191]};
    
    wire lut_1627_out = lut_1627_table[lut_1627_select];
    
    generate
    if ( USE_REG ) begin : ff_1627
        reg   lut_1627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1627_ff <= lut_1627_out;
            end
        end
        
        assign out_data[1627] = lut_1627_ff;
    end
    else begin : no_ff_1627
        assign out_data[1627] = lut_1627_out;
    end
    endgenerate
    
    
    
    // LUT : 1628
    wire [63:0] lut_1628_table = 64'b0000000000000000000000110011001100000000000000000000001110110011;
    wire [5:0] lut_1628_select = {
                             in_data[144],
                             in_data[176],
                             in_data[569],
                             in_data[543],
                             in_data[550],
                             in_data[394]};
    
    wire lut_1628_out = lut_1628_table[lut_1628_select];
    
    generate
    if ( USE_REG ) begin : ff_1628
        reg   lut_1628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1628_ff <= lut_1628_out;
            end
        end
        
        assign out_data[1628] = lut_1628_ff;
    end
    else begin : no_ff_1628
        assign out_data[1628] = lut_1628_out;
    end
    endgenerate
    
    
    
    // LUT : 1629
    wire [63:0] lut_1629_table = 64'b0000000011111111010000001111111100000000111111111100000011111111;
    wire [5:0] lut_1629_select = {
                             in_data[334],
                             in_data[488],
                             in_data[464],
                             in_data[445],
                             in_data[643],
                             in_data[732]};
    
    wire lut_1629_out = lut_1629_table[lut_1629_select];
    
    generate
    if ( USE_REG ) begin : ff_1629
        reg   lut_1629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1629_ff <= lut_1629_out;
            end
        end
        
        assign out_data[1629] = lut_1629_ff;
    end
    else begin : no_ff_1629
        assign out_data[1629] = lut_1629_out;
    end
    endgenerate
    
    
    
    // LUT : 1630
    wire [63:0] lut_1630_table = 64'b1111111100001101111111110000110111111111000000001111111100000000;
    wire [5:0] lut_1630_select = {
                             in_data[613],
                             in_data[703],
                             in_data[425],
                             in_data[718],
                             in_data[365],
                             in_data[260]};
    
    wire lut_1630_out = lut_1630_table[lut_1630_select];
    
    generate
    if ( USE_REG ) begin : ff_1630
        reg   lut_1630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1630_ff <= lut_1630_out;
            end
        end
        
        assign out_data[1630] = lut_1630_ff;
    end
    else begin : no_ff_1630
        assign out_data[1630] = lut_1630_out;
    end
    endgenerate
    
    
    
    // LUT : 1631
    wire [63:0] lut_1631_table = 64'b0000000010101011000000001010101100000000101110110000000010111011;
    wire [5:0] lut_1631_select = {
                             in_data[42],
                             in_data[139],
                             in_data[466],
                             in_data[117],
                             in_data[529],
                             in_data[546]};
    
    wire lut_1631_out = lut_1631_table[lut_1631_select];
    
    generate
    if ( USE_REG ) begin : ff_1631
        reg   lut_1631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1631_ff <= lut_1631_out;
            end
        end
        
        assign out_data[1631] = lut_1631_ff;
    end
    else begin : no_ff_1631
        assign out_data[1631] = lut_1631_out;
    end
    endgenerate
    
    
    
    // LUT : 1632
    wire [63:0] lut_1632_table = 64'b1111111111111111111111111111000011111111111100001111111111110000;
    wire [5:0] lut_1632_select = {
                             in_data[694],
                             in_data[393],
                             in_data[607],
                             in_data[435],
                             in_data[588],
                             in_data[143]};
    
    wire lut_1632_out = lut_1632_table[lut_1632_select];
    
    generate
    if ( USE_REG ) begin : ff_1632
        reg   lut_1632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1632_ff <= lut_1632_out;
            end
        end
        
        assign out_data[1632] = lut_1632_ff;
    end
    else begin : no_ff_1632
        assign out_data[1632] = lut_1632_out;
    end
    endgenerate
    
    
    
    // LUT : 1633
    wire [63:0] lut_1633_table = 64'b1110111111111111111111111111111011001111111111111100111110001100;
    wire [5:0] lut_1633_select = {
                             in_data[514],
                             in_data[522],
                             in_data[180],
                             in_data[300],
                             in_data[666],
                             in_data[368]};
    
    wire lut_1633_out = lut_1633_table[lut_1633_select];
    
    generate
    if ( USE_REG ) begin : ff_1633
        reg   lut_1633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1633_ff <= lut_1633_out;
            end
        end
        
        assign out_data[1633] = lut_1633_ff;
    end
    else begin : no_ff_1633
        assign out_data[1633] = lut_1633_out;
    end
    endgenerate
    
    
    
    // LUT : 1634
    wire [63:0] lut_1634_table = 64'b1110111111111111000000000000000011111111111111110000000011111111;
    wire [5:0] lut_1634_select = {
                             in_data[451],
                             in_data[427],
                             in_data[548],
                             in_data[309],
                             in_data[7],
                             in_data[92]};
    
    wire lut_1634_out = lut_1634_table[lut_1634_select];
    
    generate
    if ( USE_REG ) begin : ff_1634
        reg   lut_1634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1634_ff <= lut_1634_out;
            end
        end
        
        assign out_data[1634] = lut_1634_ff;
    end
    else begin : no_ff_1634
        assign out_data[1634] = lut_1634_out;
    end
    endgenerate
    
    
    
    // LUT : 1635
    wire [63:0] lut_1635_table = 64'b0000000000000000000000000000000011110011000000001111111100000000;
    wire [5:0] lut_1635_select = {
                             in_data[712],
                             in_data[649],
                             in_data[352],
                             in_data[436],
                             in_data[604],
                             in_data[639]};
    
    wire lut_1635_out = lut_1635_table[lut_1635_select];
    
    generate
    if ( USE_REG ) begin : ff_1635
        reg   lut_1635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1635_ff <= lut_1635_out;
            end
        end
        
        assign out_data[1635] = lut_1635_ff;
    end
    else begin : no_ff_1635
        assign out_data[1635] = lut_1635_out;
    end
    endgenerate
    
    
    
    // LUT : 1636
    wire [63:0] lut_1636_table = 64'b1111111111001100111111111111111111111111000000001111111111111111;
    wire [5:0] lut_1636_select = {
                             in_data[133],
                             in_data[242],
                             in_data[555],
                             in_data[762],
                             in_data[73],
                             in_data[279]};
    
    wire lut_1636_out = lut_1636_table[lut_1636_select];
    
    generate
    if ( USE_REG ) begin : ff_1636
        reg   lut_1636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1636_ff <= lut_1636_out;
            end
        end
        
        assign out_data[1636] = lut_1636_ff;
    end
    else begin : no_ff_1636
        assign out_data[1636] = lut_1636_out;
    end
    endgenerate
    
    
    
    // LUT : 1637
    wire [63:0] lut_1637_table = 64'b1111111111111111111000001111000011111111111111111111111111111111;
    wire [5:0] lut_1637_select = {
                             in_data[455],
                             in_data[304],
                             in_data[374],
                             in_data[716],
                             in_data[695],
                             in_data[371]};
    
    wire lut_1637_out = lut_1637_table[lut_1637_select];
    
    generate
    if ( USE_REG ) begin : ff_1637
        reg   lut_1637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1637_ff <= lut_1637_out;
            end
        end
        
        assign out_data[1637] = lut_1637_ff;
    end
    else begin : no_ff_1637
        assign out_data[1637] = lut_1637_out;
    end
    endgenerate
    
    
    
    // LUT : 1638
    wire [63:0] lut_1638_table = 64'b0000111001010111000010100001011100011111000101110001101100010011;
    wire [5:0] lut_1638_select = {
                             in_data[132],
                             in_data[742],
                             in_data[580],
                             in_data[452],
                             in_data[437],
                             in_data[518]};
    
    wire lut_1638_out = lut_1638_table[lut_1638_select];
    
    generate
    if ( USE_REG ) begin : ff_1638
        reg   lut_1638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1638_ff <= lut_1638_out;
            end
        end
        
        assign out_data[1638] = lut_1638_ff;
    end
    else begin : no_ff_1638
        assign out_data[1638] = lut_1638_out;
    end
    endgenerate
    
    
    
    // LUT : 1639
    wire [63:0] lut_1639_table = 64'b0000000000110000111111111111000000000001001101001111111111110100;
    wire [5:0] lut_1639_select = {
                             in_data[302],
                             in_data[605],
                             in_data[634],
                             in_data[377],
                             in_data[130],
                             in_data[775]};
    
    wire lut_1639_out = lut_1639_table[lut_1639_select];
    
    generate
    if ( USE_REG ) begin : ff_1639
        reg   lut_1639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1639_ff <= lut_1639_out;
            end
        end
        
        assign out_data[1639] = lut_1639_ff;
    end
    else begin : no_ff_1639
        assign out_data[1639] = lut_1639_out;
    end
    endgenerate
    
    
    
    // LUT : 1640
    wire [63:0] lut_1640_table = 64'b1110111011101110110011101110110011101110111011101110111011101100;
    wire [5:0] lut_1640_select = {
                             in_data[731],
                             in_data[312],
                             in_data[49],
                             in_data[673],
                             in_data[270],
                             in_data[353]};
    
    wire lut_1640_out = lut_1640_table[lut_1640_select];
    
    generate
    if ( USE_REG ) begin : ff_1640
        reg   lut_1640_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1640_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1640_ff <= lut_1640_out;
            end
        end
        
        assign out_data[1640] = lut_1640_ff;
    end
    else begin : no_ff_1640
        assign out_data[1640] = lut_1640_out;
    end
    endgenerate
    
    
    
    // LUT : 1641
    wire [63:0] lut_1641_table = 64'b1110111011101110111011101110111011101110111011101110111011101110;
    wire [5:0] lut_1641_select = {
                             in_data[142],
                             in_data[344],
                             in_data[447],
                             in_data[40],
                             in_data[630],
                             in_data[581]};
    
    wire lut_1641_out = lut_1641_table[lut_1641_select];
    
    generate
    if ( USE_REG ) begin : ff_1641
        reg   lut_1641_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1641_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1641_ff <= lut_1641_out;
            end
        end
        
        assign out_data[1641] = lut_1641_ff;
    end
    else begin : no_ff_1641
        assign out_data[1641] = lut_1641_out;
    end
    endgenerate
    
    
    
    // LUT : 1642
    wire [63:0] lut_1642_table = 64'b0000011100000111000000000000000000000111000001110000011100000111;
    wire [5:0] lut_1642_select = {
                             in_data[595],
                             in_data[583],
                             in_data[199],
                             in_data[188],
                             in_data[641],
                             in_data[370]};
    
    wire lut_1642_out = lut_1642_table[lut_1642_select];
    
    generate
    if ( USE_REG ) begin : ff_1642
        reg   lut_1642_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1642_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1642_ff <= lut_1642_out;
            end
        end
        
        assign out_data[1642] = lut_1642_ff;
    end
    else begin : no_ff_1642
        assign out_data[1642] = lut_1642_out;
    end
    endgenerate
    
    
    
    // LUT : 1643
    wire [63:0] lut_1643_table = 64'b0000111100001111000011000000110011111111111111111100111111001111;
    wire [5:0] lut_1643_select = {
                             in_data[285],
                             in_data[127],
                             in_data[278],
                             in_data[317],
                             in_data[498],
                             in_data[198]};
    
    wire lut_1643_out = lut_1643_table[lut_1643_select];
    
    generate
    if ( USE_REG ) begin : ff_1643
        reg   lut_1643_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1643_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1643_ff <= lut_1643_out;
            end
        end
        
        assign out_data[1643] = lut_1643_ff;
    end
    else begin : no_ff_1643
        assign out_data[1643] = lut_1643_out;
    end
    endgenerate
    
    
    
    // LUT : 1644
    wire [63:0] lut_1644_table = 64'b0101010101010101010101010001010101010101010101010101010100010101;
    wire [5:0] lut_1644_select = {
                             in_data[53],
                             in_data[748],
                             in_data[289],
                             in_data[307],
                             in_data[81],
                             in_data[271]};
    
    wire lut_1644_out = lut_1644_table[lut_1644_select];
    
    generate
    if ( USE_REG ) begin : ff_1644
        reg   lut_1644_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1644_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1644_ff <= lut_1644_out;
            end
        end
        
        assign out_data[1644] = lut_1644_ff;
    end
    else begin : no_ff_1644
        assign out_data[1644] = lut_1644_out;
    end
    endgenerate
    
    
    
    // LUT : 1645
    wire [63:0] lut_1645_table = 64'b1111100000001110001100000000111011111010101111111011000000111111;
    wire [5:0] lut_1645_select = {
                             in_data[174],
                             in_data[379],
                             in_data[124],
                             in_data[263],
                             in_data[491],
                             in_data[163]};
    
    wire lut_1645_out = lut_1645_table[lut_1645_select];
    
    generate
    if ( USE_REG ) begin : ff_1645
        reg   lut_1645_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1645_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1645_ff <= lut_1645_out;
            end
        end
        
        assign out_data[1645] = lut_1645_ff;
    end
    else begin : no_ff_1645
        assign out_data[1645] = lut_1645_out;
    end
    endgenerate
    
    
    
    // LUT : 1646
    wire [63:0] lut_1646_table = 64'b0001000000010000010100000101000000010000000100000101000001010000;
    wire [5:0] lut_1646_select = {
                             in_data[778],
                             in_data[72],
                             in_data[89],
                             in_data[237],
                             in_data[553],
                             in_data[178]};
    
    wire lut_1646_out = lut_1646_table[lut_1646_select];
    
    generate
    if ( USE_REG ) begin : ff_1646
        reg   lut_1646_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1646_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1646_ff <= lut_1646_out;
            end
        end
        
        assign out_data[1646] = lut_1646_ff;
    end
    else begin : no_ff_1646
        assign out_data[1646] = lut_1646_out;
    end
    endgenerate
    
    
    
    // LUT : 1647
    wire [63:0] lut_1647_table = 64'b1111111111111111111111111111111100000000000011000000110011001100;
    wire [5:0] lut_1647_select = {
                             in_data[489],
                             in_data[480],
                             in_data[120],
                             in_data[656],
                             in_data[104],
                             in_data[610]};
    
    wire lut_1647_out = lut_1647_table[lut_1647_select];
    
    generate
    if ( USE_REG ) begin : ff_1647
        reg   lut_1647_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1647_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1647_ff <= lut_1647_out;
            end
        end
        
        assign out_data[1647] = lut_1647_ff;
    end
    else begin : no_ff_1647
        assign out_data[1647] = lut_1647_out;
    end
    endgenerate
    
    
    
    // LUT : 1648
    wire [63:0] lut_1648_table = 64'b1010101000000010101010100000101010101010000000101010101000001010;
    wire [5:0] lut_1648_select = {
                             in_data[36],
                             in_data[254],
                             in_data[511],
                             in_data[592],
                             in_data[771],
                             in_data[407]};
    
    wire lut_1648_out = lut_1648_table[lut_1648_select];
    
    generate
    if ( USE_REG ) begin : ff_1648
        reg   lut_1648_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1648_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1648_ff <= lut_1648_out;
            end
        end
        
        assign out_data[1648] = lut_1648_ff;
    end
    else begin : no_ff_1648
        assign out_data[1648] = lut_1648_out;
    end
    endgenerate
    
    
    
    // LUT : 1649
    wire [63:0] lut_1649_table = 64'b1111111111111111110000001100000011111101111111111111110011111100;
    wire [5:0] lut_1649_select = {
                             in_data[651],
                             in_data[155],
                             in_data[422],
                             in_data[507],
                             in_data[501],
                             in_data[384]};
    
    wire lut_1649_out = lut_1649_table[lut_1649_select];
    
    generate
    if ( USE_REG ) begin : ff_1649
        reg   lut_1649_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1649_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1649_ff <= lut_1649_out;
            end
        end
        
        assign out_data[1649] = lut_1649_ff;
    end
    else begin : no_ff_1649
        assign out_data[1649] = lut_1649_out;
    end
    endgenerate
    
    
    
    // LUT : 1650
    wire [63:0] lut_1650_table = 64'b0101000000000000010100000001000011110001011100001111000101110001;
    wire [5:0] lut_1650_select = {
                             in_data[388],
                             in_data[310],
                             in_data[654],
                             in_data[247],
                             in_data[204],
                             in_data[96]};
    
    wire lut_1650_out = lut_1650_table[lut_1650_select];
    
    generate
    if ( USE_REG ) begin : ff_1650
        reg   lut_1650_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1650_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1650_ff <= lut_1650_out;
            end
        end
        
        assign out_data[1650] = lut_1650_ff;
    end
    else begin : no_ff_1650
        assign out_data[1650] = lut_1650_out;
    end
    endgenerate
    
    
    
    // LUT : 1651
    wire [63:0] lut_1651_table = 64'b0000111100111111000011110011111100000000000000110000000000000011;
    wire [5:0] lut_1651_select = {
                             in_data[743],
                             in_data[338],
                             in_data[454],
                             in_data[100],
                             in_data[627],
                             in_data[11]};
    
    wire lut_1651_out = lut_1651_table[lut_1651_select];
    
    generate
    if ( USE_REG ) begin : ff_1651
        reg   lut_1651_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1651_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1651_ff <= lut_1651_out;
            end
        end
        
        assign out_data[1651] = lut_1651_ff;
    end
    else begin : no_ff_1651
        assign out_data[1651] = lut_1651_out;
    end
    endgenerate
    
    
    
    // LUT : 1652
    wire [63:0] lut_1652_table = 64'b0000000000000011000000000000000000000000001100110000000000110011;
    wire [5:0] lut_1652_select = {
                             in_data[628],
                             in_data[161],
                             in_data[563],
                             in_data[184],
                             in_data[305],
                             in_data[560]};
    
    wire lut_1652_out = lut_1652_table[lut_1652_select];
    
    generate
    if ( USE_REG ) begin : ff_1652
        reg   lut_1652_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1652_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1652_ff <= lut_1652_out;
            end
        end
        
        assign out_data[1652] = lut_1652_ff;
    end
    else begin : no_ff_1652
        assign out_data[1652] = lut_1652_out;
    end
    endgenerate
    
    
    
    // LUT : 1653
    wire [63:0] lut_1653_table = 64'b0000000000000000000000001010011100000000000000000000000011110111;
    wire [5:0] lut_1653_select = {
                             in_data[670],
                             in_data[129],
                             in_data[622],
                             in_data[109],
                             in_data[38],
                             in_data[781]};
    
    wire lut_1653_out = lut_1653_table[lut_1653_select];
    
    generate
    if ( USE_REG ) begin : ff_1653
        reg   lut_1653_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1653_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1653_ff <= lut_1653_out;
            end
        end
        
        assign out_data[1653] = lut_1653_ff;
    end
    else begin : no_ff_1653
        assign out_data[1653] = lut_1653_out;
    end
    endgenerate
    
    
    
    // LUT : 1654
    wire [63:0] lut_1654_table = 64'b1100110111011101110011011101110111001100110111011100110011011101;
    wire [5:0] lut_1654_select = {
                             in_data[367],
                             in_data[674],
                             in_data[408],
                             in_data[638],
                             in_data[386],
                             in_data[152]};
    
    wire lut_1654_out = lut_1654_table[lut_1654_select];
    
    generate
    if ( USE_REG ) begin : ff_1654
        reg   lut_1654_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1654_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1654_ff <= lut_1654_out;
            end
        end
        
        assign out_data[1654] = lut_1654_ff;
    end
    else begin : no_ff_1654
        assign out_data[1654] = lut_1654_out;
    end
    endgenerate
    
    
    
    // LUT : 1655
    wire [63:0] lut_1655_table = 64'b0011001100110011101100110011001100110011001100110111001100110011;
    wire [5:0] lut_1655_select = {
                             in_data[556],
                             in_data[586],
                             in_data[125],
                             in_data[568],
                             in_data[513],
                             in_data[391]};
    
    wire lut_1655_out = lut_1655_table[lut_1655_select];
    
    generate
    if ( USE_REG ) begin : ff_1655
        reg   lut_1655_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1655_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1655_ff <= lut_1655_out;
            end
        end
        
        assign out_data[1655] = lut_1655_ff;
    end
    else begin : no_ff_1655
        assign out_data[1655] = lut_1655_out;
    end
    endgenerate
    
    
    
    // LUT : 1656
    wire [63:0] lut_1656_table = 64'b1111111111111111000011001000110000001010111111110000000000000100;
    wire [5:0] lut_1656_select = {
                             in_data[707],
                             in_data[515],
                             in_data[359],
                             in_data[43],
                             in_data[354],
                             in_data[779]};
    
    wire lut_1656_out = lut_1656_table[lut_1656_select];
    
    generate
    if ( USE_REG ) begin : ff_1656
        reg   lut_1656_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1656_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1656_ff <= lut_1656_out;
            end
        end
        
        assign out_data[1656] = lut_1656_ff;
    end
    else begin : no_ff_1656
        assign out_data[1656] = lut_1656_out;
    end
    endgenerate
    
    
    
    // LUT : 1657
    wire [63:0] lut_1657_table = 64'b0000111110001111000000000000000010001111110111110000000000000000;
    wire [5:0] lut_1657_select = {
                             in_data[118],
                             in_data[655],
                             in_data[360],
                             in_data[232],
                             in_data[539],
                             in_data[8]};
    
    wire lut_1657_out = lut_1657_table[lut_1657_select];
    
    generate
    if ( USE_REG ) begin : ff_1657
        reg   lut_1657_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1657_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1657_ff <= lut_1657_out;
            end
        end
        
        assign out_data[1657] = lut_1657_ff;
    end
    else begin : no_ff_1657
        assign out_data[1657] = lut_1657_out;
    end
    endgenerate
    
    
    
    // LUT : 1658
    wire [63:0] lut_1658_table = 64'b0101000101010001010100000101000101010001010100010101000001010001;
    wire [5:0] lut_1658_select = {
                             in_data[753],
                             in_data[726],
                             in_data[22],
                             in_data[396],
                             in_data[274],
                             in_data[122]};
    
    wire lut_1658_out = lut_1658_table[lut_1658_select];
    
    generate
    if ( USE_REG ) begin : ff_1658
        reg   lut_1658_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1658_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1658_ff <= lut_1658_out;
            end
        end
        
        assign out_data[1658] = lut_1658_ff;
    end
    else begin : no_ff_1658
        assign out_data[1658] = lut_1658_out;
    end
    endgenerate
    
    
    
    // LUT : 1659
    wire [63:0] lut_1659_table = 64'b1010101011110010000000001111000100000000111111110000000011111111;
    wire [5:0] lut_1659_select = {
                             in_data[463],
                             in_data[527],
                             in_data[290],
                             in_data[229],
                             in_data[531],
                             in_data[438]};
    
    wire lut_1659_out = lut_1659_table[lut_1659_select];
    
    generate
    if ( USE_REG ) begin : ff_1659
        reg   lut_1659_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1659_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1659_ff <= lut_1659_out;
            end
        end
        
        assign out_data[1659] = lut_1659_ff;
    end
    else begin : no_ff_1659
        assign out_data[1659] = lut_1659_out;
    end
    endgenerate
    
    
    
    // LUT : 1660
    wire [63:0] lut_1660_table = 64'b1111111111111111111111111111111111011100110111011101110011011101;
    wire [5:0] lut_1660_select = {
                             in_data[164],
                             in_data[47],
                             in_data[65],
                             in_data[534],
                             in_data[173],
                             in_data[426]};
    
    wire lut_1660_out = lut_1660_table[lut_1660_select];
    
    generate
    if ( USE_REG ) begin : ff_1660
        reg   lut_1660_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1660_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1660_ff <= lut_1660_out;
            end
        end
        
        assign out_data[1660] = lut_1660_ff;
    end
    else begin : no_ff_1660
        assign out_data[1660] = lut_1660_out;
    end
    endgenerate
    
    
    
    // LUT : 1661
    wire [63:0] lut_1661_table = 64'b0100000000000000010101010000000101000101000000000111011101000111;
    wire [5:0] lut_1661_select = {
                             in_data[720],
                             in_data[459],
                             in_data[650],
                             in_data[460],
                             in_data[154],
                             in_data[303]};
    
    wire lut_1661_out = lut_1661_table[lut_1661_select];
    
    generate
    if ( USE_REG ) begin : ff_1661
        reg   lut_1661_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1661_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1661_ff <= lut_1661_out;
            end
        end
        
        assign out_data[1661] = lut_1661_ff;
    end
    else begin : no_ff_1661
        assign out_data[1661] = lut_1661_out;
    end
    endgenerate
    
    
    
    // LUT : 1662
    wire [63:0] lut_1662_table = 64'b0000000000000000000000001000110000000000100010000000000011111111;
    wire [5:0] lut_1662_select = {
                             in_data[149],
                             in_data[283],
                             in_data[286],
                             in_data[86],
                             in_data[424],
                             in_data[67]};
    
    wire lut_1662_out = lut_1662_table[lut_1662_select];
    
    generate
    if ( USE_REG ) begin : ff_1662
        reg   lut_1662_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1662_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1662_ff <= lut_1662_out;
            end
        end
        
        assign out_data[1662] = lut_1662_ff;
    end
    else begin : no_ff_1662
        assign out_data[1662] = lut_1662_out;
    end
    endgenerate
    
    
    
    // LUT : 1663
    wire [63:0] lut_1663_table = 64'b1100110011111111000000000011001100000000110011000000000000000000;
    wire [5:0] lut_1663_select = {
                             in_data[536],
                             in_data[493],
                             in_data[710],
                             in_data[10],
                             in_data[410],
                             in_data[669]};
    
    wire lut_1663_out = lut_1663_table[lut_1663_select];
    
    generate
    if ( USE_REG ) begin : ff_1663
        reg   lut_1663_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1663_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1663_ff <= lut_1663_out;
            end
        end
        
        assign out_data[1663] = lut_1663_ff;
    end
    else begin : no_ff_1663
        assign out_data[1663] = lut_1663_out;
    end
    endgenerate
    
    
    
    // LUT : 1664
    wire [63:0] lut_1664_table = 64'b0000000010101110000000001111111100000000101011100000000011111111;
    wire [5:0] lut_1664_select = {
                             in_data[618],
                             in_data[269],
                             in_data[293],
                             in_data[147],
                             in_data[136],
                             in_data[203]};
    
    wire lut_1664_out = lut_1664_table[lut_1664_select];
    
    generate
    if ( USE_REG ) begin : ff_1664
        reg   lut_1664_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1664_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1664_ff <= lut_1664_out;
            end
        end
        
        assign out_data[1664] = lut_1664_ff;
    end
    else begin : no_ff_1664
        assign out_data[1664] = lut_1664_out;
    end
    endgenerate
    
    
    
    // LUT : 1665
    wire [63:0] lut_1665_table = 64'b0010001000110011001000100011001100100010001100110011001100110011;
    wire [5:0] lut_1665_select = {
                             in_data[168],
                             in_data[5],
                             in_data[567],
                             in_data[13],
                             in_data[351],
                             in_data[78]};
    
    wire lut_1665_out = lut_1665_table[lut_1665_select];
    
    generate
    if ( USE_REG ) begin : ff_1665
        reg   lut_1665_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1665_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1665_ff <= lut_1665_out;
            end
        end
        
        assign out_data[1665] = lut_1665_ff;
    end
    else begin : no_ff_1665
        assign out_data[1665] = lut_1665_out;
    end
    endgenerate
    
    
    
    // LUT : 1666
    wire [63:0] lut_1666_table = 64'b0000000000001100000000000000000011111111111111110000110011111111;
    wire [5:0] lut_1666_select = {
                             in_data[378],
                             in_data[159],
                             in_data[738],
                             in_data[475],
                             in_data[721],
                             in_data[29]};
    
    wire lut_1666_out = lut_1666_table[lut_1666_select];
    
    generate
    if ( USE_REG ) begin : ff_1666
        reg   lut_1666_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1666_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1666_ff <= lut_1666_out;
            end
        end
        
        assign out_data[1666] = lut_1666_ff;
    end
    else begin : no_ff_1666
        assign out_data[1666] = lut_1666_out;
    end
    endgenerate
    
    
    
    // LUT : 1667
    wire [63:0] lut_1667_table = 64'b1010111111101111000011000000110010001110110011111000110010001100;
    wire [5:0] lut_1667_select = {
                             in_data[261],
                             in_data[609],
                             in_data[416],
                             in_data[540],
                             in_data[181],
                             in_data[256]};
    
    wire lut_1667_out = lut_1667_table[lut_1667_select];
    
    generate
    if ( USE_REG ) begin : ff_1667
        reg   lut_1667_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1667_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1667_ff <= lut_1667_out;
            end
        end
        
        assign out_data[1667] = lut_1667_ff;
    end
    else begin : no_ff_1667
        assign out_data[1667] = lut_1667_out;
    end
    endgenerate
    
    
    
    // LUT : 1668
    wire [63:0] lut_1668_table = 64'b0000000000000000000000100000001000000000000000000000001000001011;
    wire [5:0] lut_1668_select = {
                             in_data[736],
                             in_data[276],
                             in_data[692],
                             in_data[244],
                             in_data[301],
                             in_data[387]};
    
    wire lut_1668_out = lut_1668_table[lut_1668_select];
    
    generate
    if ( USE_REG ) begin : ff_1668
        reg   lut_1668_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1668_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1668_ff <= lut_1668_out;
            end
        end
        
        assign out_data[1668] = lut_1668_ff;
    end
    else begin : no_ff_1668
        assign out_data[1668] = lut_1668_out;
    end
    endgenerate
    
    
    
    // LUT : 1669
    wire [63:0] lut_1669_table = 64'b1010101010001000000000000000000011111111111111111111111110111111;
    wire [5:0] lut_1669_select = {
                             in_data[443],
                             in_data[221],
                             in_data[735],
                             in_data[140],
                             in_data[380],
                             in_data[737]};
    
    wire lut_1669_out = lut_1669_table[lut_1669_select];
    
    generate
    if ( USE_REG ) begin : ff_1669
        reg   lut_1669_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1669_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1669_ff <= lut_1669_out;
            end
        end
        
        assign out_data[1669] = lut_1669_ff;
    end
    else begin : no_ff_1669
        assign out_data[1669] = lut_1669_out;
    end
    endgenerate
    
    
    
    // LUT : 1670
    wire [63:0] lut_1670_table = 64'b1111111111111111111101111111111101110111011101110100010001010101;
    wire [5:0] lut_1670_select = {
                             in_data[715],
                             in_data[70],
                             in_data[227],
                             in_data[478],
                             in_data[663],
                             in_data[494]};
    
    wire lut_1670_out = lut_1670_table[lut_1670_select];
    
    generate
    if ( USE_REG ) begin : ff_1670
        reg   lut_1670_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1670_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1670_ff <= lut_1670_out;
            end
        end
        
        assign out_data[1670] = lut_1670_ff;
    end
    else begin : no_ff_1670
        assign out_data[1670] = lut_1670_out;
    end
    endgenerate
    
    
    
    // LUT : 1671
    wire [63:0] lut_1671_table = 64'b1100110011111100110011001111110011111111111111111111111111111111;
    wire [5:0] lut_1671_select = {
                             in_data[409],
                             in_data[4],
                             in_data[606],
                             in_data[648],
                             in_data[682],
                             in_data[761]};
    
    wire lut_1671_out = lut_1671_table[lut_1671_select];
    
    generate
    if ( USE_REG ) begin : ff_1671
        reg   lut_1671_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1671_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1671_ff <= lut_1671_out;
            end
        end
        
        assign out_data[1671] = lut_1671_ff;
    end
    else begin : no_ff_1671
        assign out_data[1671] = lut_1671_out;
    end
    endgenerate
    
    
    
    // LUT : 1672
    wire [63:0] lut_1672_table = 64'b0000000000000000001000010000000000000000000000000000000100000000;
    wire [5:0] lut_1672_select = {
                             in_data[615],
                             in_data[766],
                             in_data[169],
                             in_data[33],
                             in_data[332],
                             in_data[14]};
    
    wire lut_1672_out = lut_1672_table[lut_1672_select];
    
    generate
    if ( USE_REG ) begin : ff_1672
        reg   lut_1672_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1672_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1672_ff <= lut_1672_out;
            end
        end
        
        assign out_data[1672] = lut_1672_ff;
    end
    else begin : no_ff_1672
        assign out_data[1672] = lut_1672_out;
    end
    endgenerate
    
    
    
    // LUT : 1673
    wire [63:0] lut_1673_table = 64'b1111111111111111001100110011001111111111111111110011001100110011;
    wire [5:0] lut_1673_select = {
                             in_data[751],
                             in_data[291],
                             in_data[224],
                             in_data[487],
                             in_data[572],
                             in_data[395]};
    
    wire lut_1673_out = lut_1673_table[lut_1673_select];
    
    generate
    if ( USE_REG ) begin : ff_1673
        reg   lut_1673_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1673_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1673_ff <= lut_1673_out;
            end
        end
        
        assign out_data[1673] = lut_1673_ff;
    end
    else begin : no_ff_1673
        assign out_data[1673] = lut_1673_out;
    end
    endgenerate
    
    
    
    // LUT : 1674
    wire [63:0] lut_1674_table = 64'b1100110011001100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1674_select = {
                             in_data[146],
                             in_data[234],
                             in_data[366],
                             in_data[21],
                             in_data[482],
                             in_data[157]};
    
    wire lut_1674_out = lut_1674_table[lut_1674_select];
    
    generate
    if ( USE_REG ) begin : ff_1674
        reg   lut_1674_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1674_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1674_ff <= lut_1674_out;
            end
        end
        
        assign out_data[1674] = lut_1674_ff;
    end
    else begin : no_ff_1674
        assign out_data[1674] = lut_1674_out;
    end
    endgenerate
    
    
    
    // LUT : 1675
    wire [63:0] lut_1675_table = 64'b1111111111111111111111111111111111111000100000001111101010100000;
    wire [5:0] lut_1675_select = {
                             in_data[266],
                             in_data[758],
                             in_data[282],
                             in_data[267],
                             in_data[6],
                             in_data[91]};
    
    wire lut_1675_out = lut_1675_table[lut_1675_select];
    
    generate
    if ( USE_REG ) begin : ff_1675
        reg   lut_1675_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1675_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1675_ff <= lut_1675_out;
            end
        end
        
        assign out_data[1675] = lut_1675_ff;
    end
    else begin : no_ff_1675
        assign out_data[1675] = lut_1675_out;
    end
    endgenerate
    
    
    
    // LUT : 1676
    wire [63:0] lut_1676_table = 64'b0011000011110000111100001111000001110000111100000111000011110000;
    wire [5:0] lut_1676_select = {
                             in_data[57],
                             in_data[747],
                             in_data[102],
                             in_data[97],
                             in_data[250],
                             in_data[226]};
    
    wire lut_1676_out = lut_1676_table[lut_1676_select];
    
    generate
    if ( USE_REG ) begin : ff_1676
        reg   lut_1676_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1676_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1676_ff <= lut_1676_out;
            end
        end
        
        assign out_data[1676] = lut_1676_ff;
    end
    else begin : no_ff_1676
        assign out_data[1676] = lut_1676_out;
    end
    endgenerate
    
    
    
    // LUT : 1677
    wire [63:0] lut_1677_table = 64'b1111111111111111111100001111000011111111111111111111000111110000;
    wire [5:0] lut_1677_select = {
                             in_data[82],
                             in_data[189],
                             in_data[299],
                             in_data[686],
                             in_data[668],
                             in_data[765]};
    
    wire lut_1677_out = lut_1677_table[lut_1677_select];
    
    generate
    if ( USE_REG ) begin : ff_1677
        reg   lut_1677_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1677_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1677_ff <= lut_1677_out;
            end
        end
        
        assign out_data[1677] = lut_1677_ff;
    end
    else begin : no_ff_1677
        assign out_data[1677] = lut_1677_out;
    end
    endgenerate
    
    
    
    // LUT : 1678
    wire [63:0] lut_1678_table = 64'b0000101001000010001110100101001001001010010011100100101001011110;
    wire [5:0] lut_1678_select = {
                             in_data[347],
                             in_data[504],
                             in_data[349],
                             in_data[456],
                             in_data[499],
                             in_data[403]};
    
    wire lut_1678_out = lut_1678_table[lut_1678_select];
    
    generate
    if ( USE_REG ) begin : ff_1678
        reg   lut_1678_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1678_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1678_ff <= lut_1678_out;
            end
        end
        
        assign out_data[1678] = lut_1678_ff;
    end
    else begin : no_ff_1678
        assign out_data[1678] = lut_1678_out;
    end
    endgenerate
    
    
    
    // LUT : 1679
    wire [63:0] lut_1679_table = 64'b0000000001010101000000000101010100010000010101010000000001010101;
    wire [5:0] lut_1679_select = {
                             in_data[561],
                             in_data[700],
                             in_data[236],
                             in_data[335],
                             in_data[31],
                             in_data[264]};
    
    wire lut_1679_out = lut_1679_table[lut_1679_select];
    
    generate
    if ( USE_REG ) begin : ff_1679
        reg   lut_1679_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1679_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1679_ff <= lut_1679_out;
            end
        end
        
        assign out_data[1679] = lut_1679_ff;
    end
    else begin : no_ff_1679
        assign out_data[1679] = lut_1679_out;
    end
    endgenerate
    
    
    
    // LUT : 1680
    wire [63:0] lut_1680_table = 64'b1111001011111011111100101011001011110010111110101111000011110010;
    wire [5:0] lut_1680_select = {
                             in_data[421],
                             in_data[755],
                             in_data[764],
                             in_data[521],
                             in_data[750],
                             in_data[770]};
    
    wire lut_1680_out = lut_1680_table[lut_1680_select];
    
    generate
    if ( USE_REG ) begin : ff_1680
        reg   lut_1680_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1680_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1680_ff <= lut_1680_out;
            end
        end
        
        assign out_data[1680] = lut_1680_ff;
    end
    else begin : no_ff_1680
        assign out_data[1680] = lut_1680_out;
    end
    endgenerate
    
    
    
    // LUT : 1681
    wire [63:0] lut_1681_table = 64'b1110111011101010111011101110101011101111111010101110111011101010;
    wire [5:0] lut_1681_select = {
                             in_data[662],
                             in_data[587],
                             in_data[584],
                             in_data[27],
                             in_data[473],
                             in_data[486]};
    
    wire lut_1681_out = lut_1681_table[lut_1681_select];
    
    generate
    if ( USE_REG ) begin : ff_1681
        reg   lut_1681_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1681_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1681_ff <= lut_1681_out;
            end
        end
        
        assign out_data[1681] = lut_1681_ff;
    end
    else begin : no_ff_1681
        assign out_data[1681] = lut_1681_out;
    end
    endgenerate
    
    
    
    // LUT : 1682
    wire [63:0] lut_1682_table = 64'b0001000100010001000100000001000001010111010101110111001101010011;
    wire [5:0] lut_1682_select = {
                             in_data[320],
                             in_data[678],
                             in_data[196],
                             in_data[239],
                             in_data[328],
                             in_data[570]};
    
    wire lut_1682_out = lut_1682_table[lut_1682_select];
    
    generate
    if ( USE_REG ) begin : ff_1682
        reg   lut_1682_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1682_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1682_ff <= lut_1682_out;
            end
        end
        
        assign out_data[1682] = lut_1682_ff;
    end
    else begin : no_ff_1682
        assign out_data[1682] = lut_1682_out;
    end
    endgenerate
    
    
    
    // LUT : 1683
    wire [63:0] lut_1683_table = 64'b0000001100000011000000110000001100000011000000110000001100000011;
    wire [5:0] lut_1683_select = {
                             in_data[757],
                             in_data[696],
                             in_data[138],
                             in_data[245],
                             in_data[296],
                             in_data[698]};
    
    wire lut_1683_out = lut_1683_table[lut_1683_select];
    
    generate
    if ( USE_REG ) begin : ff_1683
        reg   lut_1683_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1683_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1683_ff <= lut_1683_out;
            end
        end
        
        assign out_data[1683] = lut_1683_ff;
    end
    else begin : no_ff_1683
        assign out_data[1683] = lut_1683_out;
    end
    endgenerate
    
    
    
    // LUT : 1684
    wire [63:0] lut_1684_table = 64'b0000010000000000100000001010000001010100010001001100010011010101;
    wire [5:0] lut_1684_select = {
                             in_data[321],
                             in_data[468],
                             in_data[646],
                             in_data[355],
                             in_data[434],
                             in_data[345]};
    
    wire lut_1684_out = lut_1684_table[lut_1684_select];
    
    generate
    if ( USE_REG ) begin : ff_1684
        reg   lut_1684_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1684_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1684_ff <= lut_1684_out;
            end
        end
        
        assign out_data[1684] = lut_1684_ff;
    end
    else begin : no_ff_1684
        assign out_data[1684] = lut_1684_out;
    end
    endgenerate
    
    
    
    // LUT : 1685
    wire [63:0] lut_1685_table = 64'b1111111111111111001100110000000011111111011100010011001100000000;
    wire [5:0] lut_1685_select = {
                             in_data[681],
                             in_data[209],
                             in_data[381],
                             in_data[83],
                             in_data[160],
                             in_data[756]};
    
    wire lut_1685_out = lut_1685_table[lut_1685_select];
    
    generate
    if ( USE_REG ) begin : ff_1685
        reg   lut_1685_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1685_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1685_ff <= lut_1685_out;
            end
        end
        
        assign out_data[1685] = lut_1685_ff;
    end
    else begin : no_ff_1685
        assign out_data[1685] = lut_1685_out;
    end
    endgenerate
    
    
    
    // LUT : 1686
    wire [63:0] lut_1686_table = 64'b0000000000000000000000000000000001110001111101010111000111111111;
    wire [5:0] lut_1686_select = {
                             in_data[215],
                             in_data[614],
                             in_data[566],
                             in_data[492],
                             in_data[705],
                             in_data[457]};
    
    wire lut_1686_out = lut_1686_table[lut_1686_select];
    
    generate
    if ( USE_REG ) begin : ff_1686
        reg   lut_1686_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1686_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1686_ff <= lut_1686_out;
            end
        end
        
        assign out_data[1686] = lut_1686_ff;
    end
    else begin : no_ff_1686
        assign out_data[1686] = lut_1686_out;
    end
    endgenerate
    
    
    
    // LUT : 1687
    wire [63:0] lut_1687_table = 64'b1111000011110000111100001111000011110000111100001111000011110000;
    wire [5:0] lut_1687_select = {
                             in_data[783],
                             in_data[576],
                             in_data[730],
                             in_data[512],
                             in_data[80],
                             in_data[725]};
    
    wire lut_1687_out = lut_1687_table[lut_1687_select];
    
    generate
    if ( USE_REG ) begin : ff_1687
        reg   lut_1687_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1687_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1687_ff <= lut_1687_out;
            end
        end
        
        assign out_data[1687] = lut_1687_ff;
    end
    else begin : no_ff_1687
        assign out_data[1687] = lut_1687_out;
    end
    endgenerate
    
    
    
    // LUT : 1688
    wire [63:0] lut_1688_table = 64'b0000000000000000000000000000000000001111000011110000111100001111;
    wire [5:0] lut_1688_select = {
                             in_data[103],
                             in_data[62],
                             in_data[339],
                             in_data[440],
                             in_data[772],
                             in_data[87]};
    
    wire lut_1688_out = lut_1688_table[lut_1688_select];
    
    generate
    if ( USE_REG ) begin : ff_1688
        reg   lut_1688_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1688_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1688_ff <= lut_1688_out;
            end
        end
        
        assign out_data[1688] = lut_1688_ff;
    end
    else begin : no_ff_1688
        assign out_data[1688] = lut_1688_out;
    end
    endgenerate
    
    
    
    // LUT : 1689
    wire [63:0] lut_1689_table = 64'b1100111111001111110011111101111100000000000000000000000000001100;
    wire [5:0] lut_1689_select = {
                             in_data[183],
                             in_data[107],
                             in_data[647],
                             in_data[603],
                             in_data[121],
                             in_data[701]};
    
    wire lut_1689_out = lut_1689_table[lut_1689_select];
    
    generate
    if ( USE_REG ) begin : ff_1689
        reg   lut_1689_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1689_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1689_ff <= lut_1689_out;
            end
        end
        
        assign out_data[1689] = lut_1689_ff;
    end
    else begin : no_ff_1689
        assign out_data[1689] = lut_1689_out;
    end
    endgenerate
    
    
    
    // LUT : 1690
    wire [63:0] lut_1690_table = 64'b1100110011001100110011001101110111001100110011001100110011011100;
    wire [5:0] lut_1690_select = {
                             in_data[726],
                             in_data[247],
                             in_data[665],
                             in_data[85],
                             in_data[150],
                             in_data[137]};
    
    wire lut_1690_out = lut_1690_table[lut_1690_select];
    
    generate
    if ( USE_REG ) begin : ff_1690
        reg   lut_1690_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1690_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1690_ff <= lut_1690_out;
            end
        end
        
        assign out_data[1690] = lut_1690_ff;
    end
    else begin : no_ff_1690
        assign out_data[1690] = lut_1690_out;
    end
    endgenerate
    
    
    
    // LUT : 1691
    wire [63:0] lut_1691_table = 64'b1110111011101110111111111111111110001000100010001010111010101110;
    wire [5:0] lut_1691_select = {
                             in_data[297],
                             in_data[164],
                             in_data[24],
                             in_data[514],
                             in_data[524],
                             in_data[149]};
    
    wire lut_1691_out = lut_1691_table[lut_1691_select];
    
    generate
    if ( USE_REG ) begin : ff_1691
        reg   lut_1691_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1691_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1691_ff <= lut_1691_out;
            end
        end
        
        assign out_data[1691] = lut_1691_ff;
    end
    else begin : no_ff_1691
        assign out_data[1691] = lut_1691_out;
    end
    endgenerate
    
    
    
    // LUT : 1692
    wire [63:0] lut_1692_table = 64'b0000000011111111000000000000000100000000110101010000000000000000;
    wire [5:0] lut_1692_select = {
                             in_data[382],
                             in_data[329],
                             in_data[359],
                             in_data[766],
                             in_data[9],
                             in_data[175]};
    
    wire lut_1692_out = lut_1692_table[lut_1692_select];
    
    generate
    if ( USE_REG ) begin : ff_1692
        reg   lut_1692_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1692_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1692_ff <= lut_1692_out;
            end
        end
        
        assign out_data[1692] = lut_1692_ff;
    end
    else begin : no_ff_1692
        assign out_data[1692] = lut_1692_out;
    end
    endgenerate
    
    
    
    // LUT : 1693
    wire [63:0] lut_1693_table = 64'b0100010101010101000000000100000001010101010101010000000001000001;
    wire [5:0] lut_1693_select = {
                             in_data[12],
                             in_data[688],
                             in_data[564],
                             in_data[417],
                             in_data[762],
                             in_data[608]};
    
    wire lut_1693_out = lut_1693_table[lut_1693_select];
    
    generate
    if ( USE_REG ) begin : ff_1693
        reg   lut_1693_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1693_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1693_ff <= lut_1693_out;
            end
        end
        
        assign out_data[1693] = lut_1693_ff;
    end
    else begin : no_ff_1693
        assign out_data[1693] = lut_1693_out;
    end
    endgenerate
    
    
    
    // LUT : 1694
    wire [63:0] lut_1694_table = 64'b0100010000000100000001000000000000000000000001000101010101010101;
    wire [5:0] lut_1694_select = {
                             in_data[550],
                             in_data[604],
                             in_data[672],
                             in_data[390],
                             in_data[221],
                             in_data[469]};
    
    wire lut_1694_out = lut_1694_table[lut_1694_select];
    
    generate
    if ( USE_REG ) begin : ff_1694
        reg   lut_1694_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1694_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1694_ff <= lut_1694_out;
            end
        end
        
        assign out_data[1694] = lut_1694_ff;
    end
    else begin : no_ff_1694
        assign out_data[1694] = lut_1694_out;
    end
    endgenerate
    
    
    
    // LUT : 1695
    wire [63:0] lut_1695_table = 64'b0010001000100010001000100010001000100010001000100010001000110010;
    wire [5:0] lut_1695_select = {
                             in_data[195],
                             in_data[555],
                             in_data[394],
                             in_data[697],
                             in_data[658],
                             in_data[455]};
    
    wire lut_1695_out = lut_1695_table[lut_1695_select];
    
    generate
    if ( USE_REG ) begin : ff_1695
        reg   lut_1695_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1695_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1695_ff <= lut_1695_out;
            end
        end
        
        assign out_data[1695] = lut_1695_ff;
    end
    else begin : no_ff_1695
        assign out_data[1695] = lut_1695_out;
    end
    endgenerate
    
    
    
    // LUT : 1696
    wire [63:0] lut_1696_table = 64'b1111111111111111111111111111111100001111000011110000111100001111;
    wire [5:0] lut_1696_select = {
                             in_data[219],
                             in_data[225],
                             in_data[251],
                             in_data[180],
                             in_data[502],
                             in_data[42]};
    
    wire lut_1696_out = lut_1696_table[lut_1696_select];
    
    generate
    if ( USE_REG ) begin : ff_1696
        reg   lut_1696_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1696_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1696_ff <= lut_1696_out;
            end
        end
        
        assign out_data[1696] = lut_1696_ff;
    end
    else begin : no_ff_1696
        assign out_data[1696] = lut_1696_out;
    end
    endgenerate
    
    
    
    // LUT : 1697
    wire [63:0] lut_1697_table = 64'b1111000011110000111100001111000011111011111110111111111111111010;
    wire [5:0] lut_1697_select = {
                             in_data[595],
                             in_data[505],
                             in_data[112],
                             in_data[684],
                             in_data[731],
                             in_data[31]};
    
    wire lut_1697_out = lut_1697_table[lut_1697_select];
    
    generate
    if ( USE_REG ) begin : ff_1697
        reg   lut_1697_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1697_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1697_ff <= lut_1697_out;
            end
        end
        
        assign out_data[1697] = lut_1697_ff;
    end
    else begin : no_ff_1697
        assign out_data[1697] = lut_1697_out;
    end
    endgenerate
    
    
    
    // LUT : 1698
    wire [63:0] lut_1698_table = 64'b1000110010001100000011000000110010001110100011100000111000001110;
    wire [5:0] lut_1698_select = {
                             in_data[540],
                             in_data[518],
                             in_data[647],
                             in_data[302],
                             in_data[489],
                             in_data[151]};
    
    wire lut_1698_out = lut_1698_table[lut_1698_select];
    
    generate
    if ( USE_REG ) begin : ff_1698
        reg   lut_1698_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1698_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1698_ff <= lut_1698_out;
            end
        end
        
        assign out_data[1698] = lut_1698_ff;
    end
    else begin : no_ff_1698
        assign out_data[1698] = lut_1698_out;
    end
    endgenerate
    
    
    
    // LUT : 1699
    wire [63:0] lut_1699_table = 64'b1111111111111111000010100000001001010111010111110000000000000000;
    wire [5:0] lut_1699_select = {
                             in_data[258],
                             in_data[657],
                             in_data[245],
                             in_data[107],
                             in_data[27],
                             in_data[430]};
    
    wire lut_1699_out = lut_1699_table[lut_1699_select];
    
    generate
    if ( USE_REG ) begin : ff_1699
        reg   lut_1699_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1699_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1699_ff <= lut_1699_out;
            end
        end
        
        assign out_data[1699] = lut_1699_ff;
    end
    else begin : no_ff_1699
        assign out_data[1699] = lut_1699_out;
    end
    endgenerate
    
    
    
    // LUT : 1700
    wire [63:0] lut_1700_table = 64'b1111111111111100111111111100110011111111110111001111111111111100;
    wire [5:0] lut_1700_select = {
                             in_data[422],
                             in_data[44],
                             in_data[215],
                             in_data[474],
                             in_data[227],
                             in_data[116]};
    
    wire lut_1700_out = lut_1700_table[lut_1700_select];
    
    generate
    if ( USE_REG ) begin : ff_1700
        reg   lut_1700_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1700_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1700_ff <= lut_1700_out;
            end
        end
        
        assign out_data[1700] = lut_1700_ff;
    end
    else begin : no_ff_1700
        assign out_data[1700] = lut_1700_out;
    end
    endgenerate
    
    
    
    // LUT : 1701
    wire [63:0] lut_1701_table = 64'b0010101000000000000000000000000011111010111100000000100000001010;
    wire [5:0] lut_1701_select = {
                             in_data[275],
                             in_data[406],
                             in_data[623],
                             in_data[351],
                             in_data[23],
                             in_data[132]};
    
    wire lut_1701_out = lut_1701_table[lut_1701_select];
    
    generate
    if ( USE_REG ) begin : ff_1701
        reg   lut_1701_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1701_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1701_ff <= lut_1701_out;
            end
        end
        
        assign out_data[1701] = lut_1701_ff;
    end
    else begin : no_ff_1701
        assign out_data[1701] = lut_1701_out;
    end
    endgenerate
    
    
    
    // LUT : 1702
    wire [63:0] lut_1702_table = 64'b1111110011111100111100001111110011111100111111001111000011111100;
    wire [5:0] lut_1702_select = {
                             in_data[778],
                             in_data[620],
                             in_data[704],
                             in_data[314],
                             in_data[456],
                             in_data[207]};
    
    wire lut_1702_out = lut_1702_table[lut_1702_select];
    
    generate
    if ( USE_REG ) begin : ff_1702
        reg   lut_1702_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1702_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1702_ff <= lut_1702_out;
            end
        end
        
        assign out_data[1702] = lut_1702_ff;
    end
    else begin : no_ff_1702
        assign out_data[1702] = lut_1702_out;
    end
    endgenerate
    
    
    
    // LUT : 1703
    wire [63:0] lut_1703_table = 64'b0000000000000000101010100101010100000000000000001010101001010101;
    wire [5:0] lut_1703_select = {
                             in_data[196],
                             in_data[124],
                             in_data[527],
                             in_data[38],
                             in_data[109],
                             in_data[659]};
    
    wire lut_1703_out = lut_1703_table[lut_1703_select];
    
    generate
    if ( USE_REG ) begin : ff_1703
        reg   lut_1703_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1703_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1703_ff <= lut_1703_out;
            end
        end
        
        assign out_data[1703] = lut_1703_ff;
    end
    else begin : no_ff_1703
        assign out_data[1703] = lut_1703_out;
    end
    endgenerate
    
    
    
    // LUT : 1704
    wire [63:0] lut_1704_table = 64'b0000000000000000000000000000000000000000010101010000000001010101;
    wire [5:0] lut_1704_select = {
                             in_data[103],
                             in_data[114],
                             in_data[574],
                             in_data[393],
                             in_data[21],
                             in_data[687]};
    
    wire lut_1704_out = lut_1704_table[lut_1704_select];
    
    generate
    if ( USE_REG ) begin : ff_1704
        reg   lut_1704_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1704_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1704_ff <= lut_1704_out;
            end
        end
        
        assign out_data[1704] = lut_1704_ff;
    end
    else begin : no_ff_1704
        assign out_data[1704] = lut_1704_out;
    end
    endgenerate
    
    
    
    // LUT : 1705
    wire [63:0] lut_1705_table = 64'b0000010100000101000001010000010100101111000011111010111110101111;
    wire [5:0] lut_1705_select = {
                             in_data[327],
                             in_data[55],
                             in_data[15],
                             in_data[239],
                             in_data[110],
                             in_data[321]};
    
    wire lut_1705_out = lut_1705_table[lut_1705_select];
    
    generate
    if ( USE_REG ) begin : ff_1705
        reg   lut_1705_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1705_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1705_ff <= lut_1705_out;
            end
        end
        
        assign out_data[1705] = lut_1705_ff;
    end
    else begin : no_ff_1705
        assign out_data[1705] = lut_1705_out;
    end
    endgenerate
    
    
    
    // LUT : 1706
    wire [63:0] lut_1706_table = 64'b0011001100110011001100110011001100000000001100100000000000110011;
    wire [5:0] lut_1706_select = {
                             in_data[298],
                             in_data[383],
                             in_data[557],
                             in_data[19],
                             in_data[551],
                             in_data[8]};
    
    wire lut_1706_out = lut_1706_table[lut_1706_select];
    
    generate
    if ( USE_REG ) begin : ff_1706
        reg   lut_1706_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1706_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1706_ff <= lut_1706_out;
            end
        end
        
        assign out_data[1706] = lut_1706_ff;
    end
    else begin : no_ff_1706
        assign out_data[1706] = lut_1706_out;
    end
    endgenerate
    
    
    
    // LUT : 1707
    wire [63:0] lut_1707_table = 64'b0000000001111111000100110111011100000000000001010000000000110111;
    wire [5:0] lut_1707_select = {
                             in_data[283],
                             in_data[547],
                             in_data[261],
                             in_data[613],
                             in_data[435],
                             in_data[737]};
    
    wire lut_1707_out = lut_1707_table[lut_1707_select];
    
    generate
    if ( USE_REG ) begin : ff_1707
        reg   lut_1707_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1707_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1707_ff <= lut_1707_out;
            end
        end
        
        assign out_data[1707] = lut_1707_ff;
    end
    else begin : no_ff_1707
        assign out_data[1707] = lut_1707_out;
    end
    endgenerate
    
    
    
    // LUT : 1708
    wire [63:0] lut_1708_table = 64'b1111111111111100110011001100110011111111111111111100110011001100;
    wire [5:0] lut_1708_select = {
                             in_data[263],
                             in_data[747],
                             in_data[739],
                             in_data[68],
                             in_data[345],
                             in_data[134]};
    
    wire lut_1708_out = lut_1708_table[lut_1708_select];
    
    generate
    if ( USE_REG ) begin : ff_1708
        reg   lut_1708_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1708_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1708_ff <= lut_1708_out;
            end
        end
        
        assign out_data[1708] = lut_1708_ff;
    end
    else begin : no_ff_1708
        assign out_data[1708] = lut_1708_out;
    end
    endgenerate
    
    
    
    // LUT : 1709
    wire [63:0] lut_1709_table = 64'b1111111111111111101110001111100011111110111111101111110011111100;
    wire [5:0] lut_1709_select = {
                             in_data[153],
                             in_data[667],
                             in_data[45],
                             in_data[487],
                             in_data[513],
                             in_data[634]};
    
    wire lut_1709_out = lut_1709_table[lut_1709_select];
    
    generate
    if ( USE_REG ) begin : ff_1709
        reg   lut_1709_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1709_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1709_ff <= lut_1709_out;
            end
        end
        
        assign out_data[1709] = lut_1709_ff;
    end
    else begin : no_ff_1709
        assign out_data[1709] = lut_1709_out;
    end
    endgenerate
    
    
    
    // LUT : 1710
    wire [63:0] lut_1710_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_1710_select = {
                             in_data[87],
                             in_data[259],
                             in_data[526],
                             in_data[28],
                             in_data[310],
                             in_data[702]};
    
    wire lut_1710_out = lut_1710_table[lut_1710_select];
    
    generate
    if ( USE_REG ) begin : ff_1710
        reg   lut_1710_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1710_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1710_ff <= lut_1710_out;
            end
        end
        
        assign out_data[1710] = lut_1710_ff;
    end
    else begin : no_ff_1710
        assign out_data[1710] = lut_1710_out;
    end
    endgenerate
    
    
    
    // LUT : 1711
    wire [63:0] lut_1711_table = 64'b1100110011001100111111111111111111111111111111110000111100001111;
    wire [5:0] lut_1711_select = {
                             in_data[372],
                             in_data[380],
                             in_data[755],
                             in_data[494],
                             in_data[471],
                             in_data[648]};
    
    wire lut_1711_out = lut_1711_table[lut_1711_select];
    
    generate
    if ( USE_REG ) begin : ff_1711
        reg   lut_1711_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1711_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1711_ff <= lut_1711_out;
            end
        end
        
        assign out_data[1711] = lut_1711_ff;
    end
    else begin : no_ff_1711
        assign out_data[1711] = lut_1711_out;
    end
    endgenerate
    
    
    
    // LUT : 1712
    wire [63:0] lut_1712_table = 64'b0000010101111111000001010111111100000000000100010000000000010001;
    wire [5:0] lut_1712_select = {
                             in_data[488],
                             in_data[62],
                             in_data[398],
                             in_data[183],
                             in_data[429],
                             in_data[497]};
    
    wire lut_1712_out = lut_1712_table[lut_1712_select];
    
    generate
    if ( USE_REG ) begin : ff_1712
        reg   lut_1712_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1712_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1712_ff <= lut_1712_out;
            end
        end
        
        assign out_data[1712] = lut_1712_ff;
    end
    else begin : no_ff_1712
        assign out_data[1712] = lut_1712_out;
    end
    endgenerate
    
    
    
    // LUT : 1713
    wire [63:0] lut_1713_table = 64'b1111010111110101111100001111010111110101111101011111000011110000;
    wire [5:0] lut_1713_select = {
                             in_data[533],
                             in_data[67],
                             in_data[669],
                             in_data[130],
                             in_data[725],
                             in_data[444]};
    
    wire lut_1713_out = lut_1713_table[lut_1713_select];
    
    generate
    if ( USE_REG ) begin : ff_1713
        reg   lut_1713_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1713_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1713_ff <= lut_1713_out;
            end
        end
        
        assign out_data[1713] = lut_1713_ff;
    end
    else begin : no_ff_1713
        assign out_data[1713] = lut_1713_out;
    end
    endgenerate
    
    
    
    // LUT : 1714
    wire [63:0] lut_1714_table = 64'b0100010011011101010001001101110101000100110111010100010011111101;
    wire [5:0] lut_1714_select = {
                             in_data[649],
                             in_data[53],
                             in_data[232],
                             in_data[338],
                             in_data[193],
                             in_data[352]};
    
    wire lut_1714_out = lut_1714_table[lut_1714_select];
    
    generate
    if ( USE_REG ) begin : ff_1714
        reg   lut_1714_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1714_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1714_ff <= lut_1714_out;
            end
        end
        
        assign out_data[1714] = lut_1714_ff;
    end
    else begin : no_ff_1714
        assign out_data[1714] = lut_1714_out;
    end
    endgenerate
    
    
    
    // LUT : 1715
    wire [63:0] lut_1715_table = 64'b0101010111011101010101010101010101010101110111010101010101010100;
    wire [5:0] lut_1715_select = {
                             in_data[171],
                             in_data[483],
                             in_data[437],
                             in_data[70],
                             in_data[228],
                             in_data[491]};
    
    wire lut_1715_out = lut_1715_table[lut_1715_select];
    
    generate
    if ( USE_REG ) begin : ff_1715
        reg   lut_1715_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1715_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1715_ff <= lut_1715_out;
            end
        end
        
        assign out_data[1715] = lut_1715_ff;
    end
    else begin : no_ff_1715
        assign out_data[1715] = lut_1715_out;
    end
    endgenerate
    
    
    
    // LUT : 1716
    wire [63:0] lut_1716_table = 64'b0000101000000010000010100000101000001111000011110000111100001111;
    wire [5:0] lut_1716_select = {
                             in_data[248],
                             in_data[223],
                             in_data[170],
                             in_data[326],
                             in_data[606],
                             in_data[285]};
    
    wire lut_1716_out = lut_1716_table[lut_1716_select];
    
    generate
    if ( USE_REG ) begin : ff_1716
        reg   lut_1716_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1716_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1716_ff <= lut_1716_out;
            end
        end
        
        assign out_data[1716] = lut_1716_ff;
    end
    else begin : no_ff_1716
        assign out_data[1716] = lut_1716_out;
    end
    endgenerate
    
    
    
    // LUT : 1717
    wire [63:0] lut_1717_table = 64'b0101010101010101010101010101010101010101010101010101010101010101;
    wire [5:0] lut_1717_select = {
                             in_data[775],
                             in_data[587],
                             in_data[460],
                             in_data[640],
                             in_data[238],
                             in_data[484]};
    
    wire lut_1717_out = lut_1717_table[lut_1717_select];
    
    generate
    if ( USE_REG ) begin : ff_1717
        reg   lut_1717_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1717_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1717_ff <= lut_1717_out;
            end
        end
        
        assign out_data[1717] = lut_1717_ff;
    end
    else begin : no_ff_1717
        assign out_data[1717] = lut_1717_out;
    end
    endgenerate
    
    
    
    // LUT : 1718
    wire [63:0] lut_1718_table = 64'b0000000000110011000000000011001111111111000000111111111100000011;
    wire [5:0] lut_1718_select = {
                             in_data[566],
                             in_data[756],
                             in_data[328],
                             in_data[94],
                             in_data[441],
                             in_data[475]};
    
    wire lut_1718_out = lut_1718_table[lut_1718_select];
    
    generate
    if ( USE_REG ) begin : ff_1718
        reg   lut_1718_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1718_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1718_ff <= lut_1718_out;
            end
        end
        
        assign out_data[1718] = lut_1718_ff;
    end
    else begin : no_ff_1718
        assign out_data[1718] = lut_1718_out;
    end
    endgenerate
    
    
    
    // LUT : 1719
    wire [63:0] lut_1719_table = 64'b0101010100010001010101010101000101010101000100010101010100010001;
    wire [5:0] lut_1719_select = {
                             in_data[392],
                             in_data[142],
                             in_data[148],
                             in_data[531],
                             in_data[714],
                             in_data[289]};
    
    wire lut_1719_out = lut_1719_table[lut_1719_select];
    
    generate
    if ( USE_REG ) begin : ff_1719
        reg   lut_1719_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1719_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1719_ff <= lut_1719_out;
            end
        end
        
        assign out_data[1719] = lut_1719_ff;
    end
    else begin : no_ff_1719
        assign out_data[1719] = lut_1719_out;
    end
    endgenerate
    
    
    
    // LUT : 1720
    wire [63:0] lut_1720_table = 64'b1101111100010001110111010001000111111111110111011111111111011101;
    wire [5:0] lut_1720_select = {
                             in_data[211],
                             in_data[674],
                             in_data[332],
                             in_data[37],
                             in_data[187],
                             in_data[546]};
    
    wire lut_1720_out = lut_1720_table[lut_1720_select];
    
    generate
    if ( USE_REG ) begin : ff_1720
        reg   lut_1720_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1720_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1720_ff <= lut_1720_out;
            end
        end
        
        assign out_data[1720] = lut_1720_ff;
    end
    else begin : no_ff_1720
        assign out_data[1720] = lut_1720_out;
    end
    endgenerate
    
    
    
    // LUT : 1721
    wire [63:0] lut_1721_table = 64'b1111111111111111101111111010111110101111101011111010101100101010;
    wire [5:0] lut_1721_select = {
                             in_data[173],
                             in_data[166],
                             in_data[14],
                             in_data[724],
                             in_data[92],
                             in_data[147]};
    
    wire lut_1721_out = lut_1721_table[lut_1721_select];
    
    generate
    if ( USE_REG ) begin : ff_1721
        reg   lut_1721_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1721_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1721_ff <= lut_1721_out;
            end
        end
        
        assign out_data[1721] = lut_1721_ff;
    end
    else begin : no_ff_1721
        assign out_data[1721] = lut_1721_out;
    end
    endgenerate
    
    
    
    // LUT : 1722
    wire [63:0] lut_1722_table = 64'b1010101110101011101010111010101110101011101010111010101110101011;
    wire [5:0] lut_1722_select = {
                             in_data[40],
                             in_data[5],
                             in_data[643],
                             in_data[592],
                             in_data[539],
                             in_data[161]};
    
    wire lut_1722_out = lut_1722_table[lut_1722_select];
    
    generate
    if ( USE_REG ) begin : ff_1722
        reg   lut_1722_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1722_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1722_ff <= lut_1722_out;
            end
        end
        
        assign out_data[1722] = lut_1722_ff;
    end
    else begin : no_ff_1722
        assign out_data[1722] = lut_1722_out;
    end
    endgenerate
    
    
    
    // LUT : 1723
    wire [63:0] lut_1723_table = 64'b1111111111111111101010110010001011111111101110111111101110111011;
    wire [5:0] lut_1723_select = {
                             in_data[442],
                             in_data[343],
                             in_data[230],
                             in_data[768],
                             in_data[493],
                             in_data[340]};
    
    wire lut_1723_out = lut_1723_table[lut_1723_select];
    
    generate
    if ( USE_REG ) begin : ff_1723
        reg   lut_1723_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1723_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1723_ff <= lut_1723_out;
            end
        end
        
        assign out_data[1723] = lut_1723_ff;
    end
    else begin : no_ff_1723
        assign out_data[1723] = lut_1723_out;
    end
    endgenerate
    
    
    
    // LUT : 1724
    wire [63:0] lut_1724_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_1724_select = {
                             in_data[461],
                             in_data[318],
                             in_data[288],
                             in_data[562],
                             in_data[559],
                             in_data[641]};
    
    wire lut_1724_out = lut_1724_table[lut_1724_select];
    
    generate
    if ( USE_REG ) begin : ff_1724
        reg   lut_1724_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1724_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1724_ff <= lut_1724_out;
            end
        end
        
        assign out_data[1724] = lut_1724_ff;
    end
    else begin : no_ff_1724
        assign out_data[1724] = lut_1724_out;
    end
    endgenerate
    
    
    
    // LUT : 1725
    wire [63:0] lut_1725_table = 64'b0010101100101011001000110010001000101011001110110010101100111011;
    wire [5:0] lut_1725_select = {
                             in_data[86],
                             in_data[758],
                             in_data[26],
                             in_data[303],
                             in_data[600],
                             in_data[495]};
    
    wire lut_1725_out = lut_1725_table[lut_1725_select];
    
    generate
    if ( USE_REG ) begin : ff_1725
        reg   lut_1725_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1725_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1725_ff <= lut_1725_out;
            end
        end
        
        assign out_data[1725] = lut_1725_ff;
    end
    else begin : no_ff_1725
        assign out_data[1725] = lut_1725_out;
    end
    endgenerate
    
    
    
    // LUT : 1726
    wire [63:0] lut_1726_table = 64'b1101110011111111110000001111111111000000111111111100000011111111;
    wire [5:0] lut_1726_select = {
                             in_data[1],
                             in_data[88],
                             in_data[236],
                             in_data[249],
                             in_data[736],
                             in_data[10]};
    
    wire lut_1726_out = lut_1726_table[lut_1726_select];
    
    generate
    if ( USE_REG ) begin : ff_1726
        reg   lut_1726_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1726_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1726_ff <= lut_1726_out;
            end
        end
        
        assign out_data[1726] = lut_1726_ff;
    end
    else begin : no_ff_1726
        assign out_data[1726] = lut_1726_out;
    end
    endgenerate
    
    
    
    // LUT : 1727
    wire [63:0] lut_1727_table = 64'b0011000000010000000000000000000001110111001100110000001100000011;
    wire [5:0] lut_1727_select = {
                             in_data[357],
                             in_data[74],
                             in_data[744],
                             in_data[413],
                             in_data[656],
                             in_data[91]};
    
    wire lut_1727_out = lut_1727_table[lut_1727_select];
    
    generate
    if ( USE_REG ) begin : ff_1727
        reg   lut_1727_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1727_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1727_ff <= lut_1727_out;
            end
        end
        
        assign out_data[1727] = lut_1727_ff;
    end
    else begin : no_ff_1727
        assign out_data[1727] = lut_1727_out;
    end
    endgenerate
    
    
    
    // LUT : 1728
    wire [63:0] lut_1728_table = 64'b1111001111111111001100110011001111110011111100110000000000100011;
    wire [5:0] lut_1728_select = {
                             in_data[246],
                             in_data[202],
                             in_data[580],
                             in_data[721],
                             in_data[581],
                             in_data[33]};
    
    wire lut_1728_out = lut_1728_table[lut_1728_select];
    
    generate
    if ( USE_REG ) begin : ff_1728
        reg   lut_1728_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1728_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1728_ff <= lut_1728_out;
            end
        end
        
        assign out_data[1728] = lut_1728_ff;
    end
    else begin : no_ff_1728
        assign out_data[1728] = lut_1728_out;
    end
    endgenerate
    
    
    
    // LUT : 1729
    wire [63:0] lut_1729_table = 64'b0101010100000000010101110000000011110111000000000111011100000000;
    wire [5:0] lut_1729_select = {
                             in_data[536],
                             in_data[304],
                             in_data[209],
                             in_data[397],
                             in_data[69],
                             in_data[594]};
    
    wire lut_1729_out = lut_1729_table[lut_1729_select];
    
    generate
    if ( USE_REG ) begin : ff_1729
        reg   lut_1729_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1729_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1729_ff <= lut_1729_out;
            end
        end
        
        assign out_data[1729] = lut_1729_ff;
    end
    else begin : no_ff_1729
        assign out_data[1729] = lut_1729_out;
    end
    endgenerate
    
    
    
    // LUT : 1730
    wire [63:0] lut_1730_table = 64'b1010111110101010111111111010111010101111101010101110111110101110;
    wire [5:0] lut_1730_select = {
                             in_data[560],
                             in_data[625],
                             in_data[610],
                             in_data[205],
                             in_data[186],
                             in_data[213]};
    
    wire lut_1730_out = lut_1730_table[lut_1730_select];
    
    generate
    if ( USE_REG ) begin : ff_1730
        reg   lut_1730_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1730_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1730_ff <= lut_1730_out;
            end
        end
        
        assign out_data[1730] = lut_1730_ff;
    end
    else begin : no_ff_1730
        assign out_data[1730] = lut_1730_out;
    end
    endgenerate
    
    
    
    // LUT : 1731
    wire [63:0] lut_1731_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_1731_select = {
                             in_data[676],
                             in_data[626],
                             in_data[309],
                             in_data[203],
                             in_data[750],
                             in_data[773]};
    
    wire lut_1731_out = lut_1731_table[lut_1731_select];
    
    generate
    if ( USE_REG ) begin : ff_1731
        reg   lut_1731_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1731_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1731_ff <= lut_1731_out;
            end
        end
        
        assign out_data[1731] = lut_1731_ff;
    end
    else begin : no_ff_1731
        assign out_data[1731] = lut_1731_out;
    end
    endgenerate
    
    
    
    // LUT : 1732
    wire [63:0] lut_1732_table = 64'b0010001000110011001000000011001100100000001100110000000000110011;
    wire [5:0] lut_1732_select = {
                             in_data[197],
                             in_data[671],
                             in_data[629],
                             in_data[503],
                             in_data[331],
                             in_data[389]};
    
    wire lut_1732_out = lut_1732_table[lut_1732_select];
    
    generate
    if ( USE_REG ) begin : ff_1732
        reg   lut_1732_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1732_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1732_ff <= lut_1732_out;
            end
        end
        
        assign out_data[1732] = lut_1732_ff;
    end
    else begin : no_ff_1732
        assign out_data[1732] = lut_1732_out;
    end
    endgenerate
    
    
    
    // LUT : 1733
    wire [63:0] lut_1733_table = 64'b1111111111111111011111111111111111111010111110100000000000000000;
    wire [5:0] lut_1733_select = {
                             in_data[440],
                             in_data[399],
                             in_data[507],
                             in_data[157],
                             in_data[447],
                             in_data[369]};
    
    wire lut_1733_out = lut_1733_table[lut_1733_select];
    
    generate
    if ( USE_REG ) begin : ff_1733
        reg   lut_1733_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1733_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1733_ff <= lut_1733_out;
            end
        end
        
        assign out_data[1733] = lut_1733_ff;
    end
    else begin : no_ff_1733
        assign out_data[1733] = lut_1733_out;
    end
    endgenerate
    
    
    
    // LUT : 1734
    wire [63:0] lut_1734_table = 64'b0000111100001111000011100000101000001111000011110000111100001111;
    wire [5:0] lut_1734_select = {
                             in_data[517],
                             in_data[771],
                             in_data[29],
                             in_data[685],
                             in_data[590],
                             in_data[360]};
    
    wire lut_1734_out = lut_1734_table[lut_1734_select];
    
    generate
    if ( USE_REG ) begin : ff_1734
        reg   lut_1734_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1734_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1734_ff <= lut_1734_out;
            end
        end
        
        assign out_data[1734] = lut_1734_ff;
    end
    else begin : no_ff_1734
        assign out_data[1734] = lut_1734_out;
    end
    endgenerate
    
    
    
    // LUT : 1735
    wire [63:0] lut_1735_table = 64'b0000000000000000110011001000110000000011000000110011001100111011;
    wire [5:0] lut_1735_select = {
                             in_data[409],
                             in_data[301],
                             in_data[75],
                             in_data[627],
                             in_data[519],
                             in_data[366]};
    
    wire lut_1735_out = lut_1735_table[lut_1735_select];
    
    generate
    if ( USE_REG ) begin : ff_1735
        reg   lut_1735_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1735_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1735_ff <= lut_1735_out;
            end
        end
        
        assign out_data[1735] = lut_1735_ff;
    end
    else begin : no_ff_1735
        assign out_data[1735] = lut_1735_out;
    end
    endgenerate
    
    
    
    // LUT : 1736
    wire [63:0] lut_1736_table = 64'b1110110011111101111010001111110111101111111111111100110011011101;
    wire [5:0] lut_1736_select = {
                             in_data[374],
                             in_data[633],
                             in_data[538],
                             in_data[567],
                             in_data[452],
                             in_data[354]};
    
    wire lut_1736_out = lut_1736_table[lut_1736_select];
    
    generate
    if ( USE_REG ) begin : ff_1736
        reg   lut_1736_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1736_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1736_ff <= lut_1736_out;
            end
        end
        
        assign out_data[1736] = lut_1736_ff;
    end
    else begin : no_ff_1736
        assign out_data[1736] = lut_1736_out;
    end
    endgenerate
    
    
    
    // LUT : 1737
    wire [63:0] lut_1737_table = 64'b0000010100000101000101110000011100000111000001010001111100000111;
    wire [5:0] lut_1737_select = {
                             in_data[138],
                             in_data[565],
                             in_data[558],
                             in_data[384],
                             in_data[772],
                             in_data[465]};
    
    wire lut_1737_out = lut_1737_table[lut_1737_select];
    
    generate
    if ( USE_REG ) begin : ff_1737
        reg   lut_1737_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1737_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1737_ff <= lut_1737_out;
            end
        end
        
        assign out_data[1737] = lut_1737_ff;
    end
    else begin : no_ff_1737
        assign out_data[1737] = lut_1737_out;
    end
    endgenerate
    
    
    
    // LUT : 1738
    wire [63:0] lut_1738_table = 64'b1111111111111111000000000001000011111111111111110000000001010000;
    wire [5:0] lut_1738_select = {
                             in_data[612],
                             in_data[182],
                             in_data[769],
                             in_data[274],
                             in_data[4],
                             in_data[25]};
    
    wire lut_1738_out = lut_1738_table[lut_1738_select];
    
    generate
    if ( USE_REG ) begin : ff_1738
        reg   lut_1738_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1738_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1738_ff <= lut_1738_out;
            end
        end
        
        assign out_data[1738] = lut_1738_ff;
    end
    else begin : no_ff_1738
        assign out_data[1738] = lut_1738_out;
    end
    endgenerate
    
    
    
    // LUT : 1739
    wire [63:0] lut_1739_table = 64'b1110111111111111000011110000111100001111111111110000000000001111;
    wire [5:0] lut_1739_select = {
                             in_data[568],
                             in_data[217],
                             in_data[233],
                             in_data[579],
                             in_data[689],
                             in_data[644]};
    
    wire lut_1739_out = lut_1739_table[lut_1739_select];
    
    generate
    if ( USE_REG ) begin : ff_1739
        reg   lut_1739_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1739_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1739_ff <= lut_1739_out;
            end
        end
        
        assign out_data[1739] = lut_1739_ff;
    end
    else begin : no_ff_1739
        assign out_data[1739] = lut_1739_out;
    end
    endgenerate
    
    
    
    // LUT : 1740
    wire [63:0] lut_1740_table = 64'b0011001100110011001100110011001100000000000000000000000000000000;
    wire [5:0] lut_1740_select = {
                             in_data[350],
                             in_data[638],
                             in_data[3],
                             in_data[499],
                             in_data[244],
                             in_data[418]};
    
    wire lut_1740_out = lut_1740_table[lut_1740_select];
    
    generate
    if ( USE_REG ) begin : ff_1740
        reg   lut_1740_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1740_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1740_ff <= lut_1740_out;
            end
        end
        
        assign out_data[1740] = lut_1740_ff;
    end
    else begin : no_ff_1740
        assign out_data[1740] = lut_1740_out;
    end
    endgenerate
    
    
    
    // LUT : 1741
    wire [63:0] lut_1741_table = 64'b1111111111111111111111111111111111110000111100101111000011110000;
    wire [5:0] lut_1741_select = {
                             in_data[152],
                             in_data[117],
                             in_data[61],
                             in_data[102],
                             in_data[458],
                             in_data[49]};
    
    wire lut_1741_out = lut_1741_table[lut_1741_select];
    
    generate
    if ( USE_REG ) begin : ff_1741
        reg   lut_1741_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1741_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1741_ff <= lut_1741_out;
            end
        end
        
        assign out_data[1741] = lut_1741_ff;
    end
    else begin : no_ff_1741
        assign out_data[1741] = lut_1741_out;
    end
    endgenerate
    
    
    
    // LUT : 1742
    wire [63:0] lut_1742_table = 64'b0101010111111111010101011111111100000000000000000000000001010101;
    wire [5:0] lut_1742_select = {
                             in_data[262],
                             in_data[424],
                             in_data[695],
                             in_data[2],
                             in_data[118],
                             in_data[570]};
    
    wire lut_1742_out = lut_1742_table[lut_1742_select];
    
    generate
    if ( USE_REG ) begin : ff_1742
        reg   lut_1742_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1742_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1742_ff <= lut_1742_out;
            end
        end
        
        assign out_data[1742] = lut_1742_ff;
    end
    else begin : no_ff_1742
        assign out_data[1742] = lut_1742_out;
    end
    endgenerate
    
    
    
    // LUT : 1743
    wire [63:0] lut_1743_table = 64'b0000000000001100000000000000110000001111000011000000111100001111;
    wire [5:0] lut_1743_select = {
                             in_data[662],
                             in_data[530],
                             in_data[463],
                             in_data[414],
                             in_data[522],
                             in_data[7]};
    
    wire lut_1743_out = lut_1743_table[lut_1743_select];
    
    generate
    if ( USE_REG ) begin : ff_1743
        reg   lut_1743_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1743_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1743_ff <= lut_1743_out;
            end
        end
        
        assign out_data[1743] = lut_1743_ff;
    end
    else begin : no_ff_1743
        assign out_data[1743] = lut_1743_out;
    end
    endgenerate
    
    
    
    // LUT : 1744
    wire [63:0] lut_1744_table = 64'b1110111011001100111111111100110011101100110011001111111111001100;
    wire [5:0] lut_1744_select = {
                             in_data[11],
                             in_data[678],
                             in_data[666],
                             in_data[602],
                             in_data[609],
                             in_data[391]};
    
    wire lut_1744_out = lut_1744_table[lut_1744_select];
    
    generate
    if ( USE_REG ) begin : ff_1744
        reg   lut_1744_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1744_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1744_ff <= lut_1744_out;
            end
        end
        
        assign out_data[1744] = lut_1744_ff;
    end
    else begin : no_ff_1744
        assign out_data[1744] = lut_1744_out;
    end
    endgenerate
    
    
    
    // LUT : 1745
    wire [63:0] lut_1745_table = 64'b0100000011110000110111011111111100000000000000001100000011110000;
    wire [5:0] lut_1745_select = {
                             in_data[273],
                             in_data[664],
                             in_data[293],
                             in_data[438],
                             in_data[325],
                             in_data[677]};
    
    wire lut_1745_out = lut_1745_table[lut_1745_select];
    
    generate
    if ( USE_REG ) begin : ff_1745
        reg   lut_1745_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1745_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1745_ff <= lut_1745_out;
            end
        end
        
        assign out_data[1745] = lut_1745_ff;
    end
    else begin : no_ff_1745
        assign out_data[1745] = lut_1745_out;
    end
    endgenerate
    
    
    
    // LUT : 1746
    wire [63:0] lut_1746_table = 64'b1100110000000000111111111111111110000100000000001111110111111111;
    wire [5:0] lut_1746_select = {
                             in_data[733],
                             in_data[408],
                             in_data[265],
                             in_data[290],
                             in_data[520],
                             in_data[556]};
    
    wire lut_1746_out = lut_1746_table[lut_1746_select];
    
    generate
    if ( USE_REG ) begin : ff_1746
        reg   lut_1746_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1746_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1746_ff <= lut_1746_out;
            end
        end
        
        assign out_data[1746] = lut_1746_ff;
    end
    else begin : no_ff_1746
        assign out_data[1746] = lut_1746_out;
    end
    endgenerate
    
    
    
    // LUT : 1747
    wire [63:0] lut_1747_table = 64'b0000111100001111000011110000111100000000000011110000000000001111;
    wire [5:0] lut_1747_select = {
                             in_data[637],
                             in_data[694],
                             in_data[267],
                             in_data[388],
                             in_data[757],
                             in_data[36]};
    
    wire lut_1747_out = lut_1747_table[lut_1747_select];
    
    generate
    if ( USE_REG ) begin : ff_1747
        reg   lut_1747_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1747_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1747_ff <= lut_1747_out;
            end
        end
        
        assign out_data[1747] = lut_1747_ff;
    end
    else begin : no_ff_1747
        assign out_data[1747] = lut_1747_out;
    end
    endgenerate
    
    
    
    // LUT : 1748
    wire [63:0] lut_1748_table = 64'b0000000011001100000000001111111100000100110011001100110011111111;
    wire [5:0] lut_1748_select = {
                             in_data[184],
                             in_data[535],
                             in_data[378],
                             in_data[333],
                             in_data[330],
                             in_data[226]};
    
    wire lut_1748_out = lut_1748_table[lut_1748_select];
    
    generate
    if ( USE_REG ) begin : ff_1748
        reg   lut_1748_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1748_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1748_ff <= lut_1748_out;
            end
        end
        
        assign out_data[1748] = lut_1748_ff;
    end
    else begin : no_ff_1748
        assign out_data[1748] = lut_1748_out;
    end
    endgenerate
    
    
    
    // LUT : 1749
    wire [63:0] lut_1749_table = 64'b1111111111111010111111111111101011111111111110101111111111111010;
    wire [5:0] lut_1749_select = {
                             in_data[361],
                             in_data[504],
                             in_data[93],
                             in_data[599],
                             in_data[252],
                             in_data[66]};
    
    wire lut_1749_out = lut_1749_table[lut_1749_select];
    
    generate
    if ( USE_REG ) begin : ff_1749
        reg   lut_1749_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1749_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1749_ff <= lut_1749_out;
            end
        end
        
        assign out_data[1749] = lut_1749_ff;
    end
    else begin : no_ff_1749
        assign out_data[1749] = lut_1749_out;
    end
    endgenerate
    
    
    
    // LUT : 1750
    wire [63:0] lut_1750_table = 64'b0000000000000000001000100010001000000000000000000010001000100010;
    wire [5:0] lut_1750_select = {
                             in_data[642],
                             in_data[194],
                             in_data[699],
                             in_data[479],
                             in_data[250],
                             in_data[515]};
    
    wire lut_1750_out = lut_1750_table[lut_1750_select];
    
    generate
    if ( USE_REG ) begin : ff_1750
        reg   lut_1750_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1750_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1750_ff <= lut_1750_out;
            end
        end
        
        assign out_data[1750] = lut_1750_ff;
    end
    else begin : no_ff_1750
        assign out_data[1750] = lut_1750_out;
    end
    endgenerate
    
    
    
    // LUT : 1751
    wire [63:0] lut_1751_table = 64'b1111111111111100111111001100000011111111111111111111111111111110;
    wire [5:0] lut_1751_select = {
                             in_data[742],
                             in_data[445],
                             in_data[621],
                             in_data[146],
                             in_data[120],
                             in_data[698]};
    
    wire lut_1751_out = lut_1751_table[lut_1751_select];
    
    generate
    if ( USE_REG ) begin : ff_1751
        reg   lut_1751_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1751_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1751_ff <= lut_1751_out;
            end
        end
        
        assign out_data[1751] = lut_1751_ff;
    end
    else begin : no_ff_1751
        assign out_data[1751] = lut_1751_out;
    end
    endgenerate
    
    
    
    // LUT : 1752
    wire [63:0] lut_1752_table = 64'b0000000000000011000000000000001100000000000011110000000000001111;
    wire [5:0] lut_1752_select = {
                             in_data[571],
                             in_data[703],
                             in_data[542],
                             in_data[190],
                             in_data[78],
                             in_data[532]};
    
    wire lut_1752_out = lut_1752_table[lut_1752_select];
    
    generate
    if ( USE_REG ) begin : ff_1752
        reg   lut_1752_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1752_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1752_ff <= lut_1752_out;
            end
        end
        
        assign out_data[1752] = lut_1752_ff;
    end
    else begin : no_ff_1752
        assign out_data[1752] = lut_1752_out;
    end
    endgenerate
    
    
    
    // LUT : 1753
    wire [63:0] lut_1753_table = 64'b1100010011110100110001001111100011000000110000001100000011111000;
    wire [5:0] lut_1753_select = {
                             in_data[201],
                             in_data[511],
                             in_data[683],
                             in_data[212],
                             in_data[601],
                             in_data[411]};
    
    wire lut_1753_out = lut_1753_table[lut_1753_select];
    
    generate
    if ( USE_REG ) begin : ff_1753
        reg   lut_1753_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1753_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1753_ff <= lut_1753_out;
            end
        end
        
        assign out_data[1753] = lut_1753_ff;
    end
    else begin : no_ff_1753
        assign out_data[1753] = lut_1753_out;
    end
    endgenerate
    
    
    
    // LUT : 1754
    wire [63:0] lut_1754_table = 64'b0000000000000000000000000000000011111110111111111111111100100010;
    wire [5:0] lut_1754_select = {
                             in_data[583],
                             in_data[428],
                             in_data[324],
                             in_data[111],
                             in_data[661],
                             in_data[423]};
    
    wire lut_1754_out = lut_1754_table[lut_1754_select];
    
    generate
    if ( USE_REG ) begin : ff_1754
        reg   lut_1754_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1754_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1754_ff <= lut_1754_out;
            end
        end
        
        assign out_data[1754] = lut_1754_ff;
    end
    else begin : no_ff_1754
        assign out_data[1754] = lut_1754_out;
    end
    endgenerate
    
    
    
    // LUT : 1755
    wire [63:0] lut_1755_table = 64'b0011001100110011001100110011001101010111000101111010101010101010;
    wire [5:0] lut_1755_select = {
                             in_data[525],
                             in_data[402],
                             in_data[473],
                             in_data[516],
                             in_data[631],
                             in_data[286]};
    
    wire lut_1755_out = lut_1755_table[lut_1755_select];
    
    generate
    if ( USE_REG ) begin : ff_1755
        reg   lut_1755_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1755_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1755_ff <= lut_1755_out;
            end
        end
        
        assign out_data[1755] = lut_1755_ff;
    end
    else begin : no_ff_1755
        assign out_data[1755] = lut_1755_out;
    end
    endgenerate
    
    
    
    // LUT : 1756
    wire [63:0] lut_1756_table = 64'b1111111011111111101110101111111110101010111111101010101010101010;
    wire [5:0] lut_1756_select = {
                             in_data[710],
                             in_data[751],
                             in_data[294],
                             in_data[81],
                             in_data[307],
                             in_data[401]};
    
    wire lut_1756_out = lut_1756_table[lut_1756_select];
    
    generate
    if ( USE_REG ) begin : ff_1756
        reg   lut_1756_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1756_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1756_ff <= lut_1756_out;
            end
        end
        
        assign out_data[1756] = lut_1756_ff;
    end
    else begin : no_ff_1756
        assign out_data[1756] = lut_1756_out;
    end
    endgenerate
    
    
    
    // LUT : 1757
    wire [63:0] lut_1757_table = 64'b0000000000000000000000000000000010101010101011101010101011101110;
    wire [5:0] lut_1757_select = {
                             in_data[257],
                             in_data[278],
                             in_data[510],
                             in_data[708],
                             in_data[572],
                             in_data[154]};
    
    wire lut_1757_out = lut_1757_table[lut_1757_select];
    
    generate
    if ( USE_REG ) begin : ff_1757
        reg   lut_1757_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1757_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1757_ff <= lut_1757_out;
            end
        end
        
        assign out_data[1757] = lut_1757_ff;
    end
    else begin : no_ff_1757
        assign out_data[1757] = lut_1757_out;
    end
    endgenerate
    
    
    
    // LUT : 1758
    wire [63:0] lut_1758_table = 64'b1111010101010000110101010101010111110101010101001111010101010101;
    wire [5:0] lut_1758_select = {
                             in_data[506],
                             in_data[191],
                             in_data[582],
                             in_data[576],
                             in_data[561],
                             in_data[158]};
    
    wire lut_1758_out = lut_1758_table[lut_1758_select];
    
    generate
    if ( USE_REG ) begin : ff_1758
        reg   lut_1758_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1758_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1758_ff <= lut_1758_out;
            end
        end
        
        assign out_data[1758] = lut_1758_ff;
    end
    else begin : no_ff_1758
        assign out_data[1758] = lut_1758_out;
    end
    endgenerate
    
    
    
    // LUT : 1759
    wire [63:0] lut_1759_table = 64'b1010101000001010010000000000000000000000000010110101000001010001;
    wire [5:0] lut_1759_select = {
                             in_data[185],
                             in_data[214],
                             in_data[549],
                             in_data[264],
                             in_data[774],
                             in_data[541]};
    
    wire lut_1759_out = lut_1759_table[lut_1759_select];
    
    generate
    if ( USE_REG ) begin : ff_1759
        reg   lut_1759_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1759_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1759_ff <= lut_1759_out;
            end
        end
        
        assign out_data[1759] = lut_1759_ff;
    end
    else begin : no_ff_1759
        assign out_data[1759] = lut_1759_out;
    end
    endgenerate
    
    
    
    // LUT : 1760
    wire [63:0] lut_1760_table = 64'b0000000000000000111111111111111100001110000011001110111011101110;
    wire [5:0] lut_1760_select = {
                             in_data[605],
                             in_data[322],
                             in_data[59],
                             in_data[554],
                             in_data[349],
                             in_data[403]};
    
    wire lut_1760_out = lut_1760_table[lut_1760_select];
    
    generate
    if ( USE_REG ) begin : ff_1760
        reg   lut_1760_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1760_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1760_ff <= lut_1760_out;
            end
        end
        
        assign out_data[1760] = lut_1760_ff;
    end
    else begin : no_ff_1760
        assign out_data[1760] = lut_1760_out;
    end
    endgenerate
    
    
    
    // LUT : 1761
    wire [63:0] lut_1761_table = 64'b0001000100010001000100110001001100010001000100010001000100010001;
    wire [5:0] lut_1761_select = {
                             in_data[6],
                             in_data[754],
                             in_data[670],
                             in_data[136],
                             in_data[268],
                             in_data[179]};
    
    wire lut_1761_out = lut_1761_table[lut_1761_select];
    
    generate
    if ( USE_REG ) begin : ff_1761
        reg   lut_1761_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1761_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1761_ff <= lut_1761_out;
            end
        end
        
        assign out_data[1761] = lut_1761_ff;
    end
    else begin : no_ff_1761
        assign out_data[1761] = lut_1761_out;
    end
    endgenerate
    
    
    
    // LUT : 1762
    wire [63:0] lut_1762_table = 64'b1111111111111111111111111111111111101110111011101010111011101110;
    wire [5:0] lut_1762_select = {
                             in_data[204],
                             in_data[614],
                             in_data[363],
                             in_data[54],
                             in_data[679],
                             in_data[121]};
    
    wire lut_1762_out = lut_1762_table[lut_1762_select];
    
    generate
    if ( USE_REG ) begin : ff_1762
        reg   lut_1762_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1762_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1762_ff <= lut_1762_out;
            end
        end
        
        assign out_data[1762] = lut_1762_ff;
    end
    else begin : no_ff_1762
        assign out_data[1762] = lut_1762_out;
    end
    endgenerate
    
    
    
    // LUT : 1763
    wire [63:0] lut_1763_table = 64'b0011001100110011000000000011001000110000001100000000000000110000;
    wire [5:0] lut_1763_select = {
                             in_data[492],
                             in_data[386],
                             in_data[611],
                             in_data[464],
                             in_data[500],
                             in_data[730]};
    
    wire lut_1763_out = lut_1763_table[lut_1763_select];
    
    generate
    if ( USE_REG ) begin : ff_1763
        reg   lut_1763_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1763_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1763_ff <= lut_1763_out;
            end
        end
        
        assign out_data[1763] = lut_1763_ff;
    end
    else begin : no_ff_1763
        assign out_data[1763] = lut_1763_out;
    end
    endgenerate
    
    
    
    // LUT : 1764
    wire [63:0] lut_1764_table = 64'b0101111100000000111111111111111111111111101000001111111111111010;
    wire [5:0] lut_1764_select = {
                             in_data[711],
                             in_data[376],
                             in_data[287],
                             in_data[260],
                             in_data[337],
                             in_data[690]};
    
    wire lut_1764_out = lut_1764_table[lut_1764_select];
    
    generate
    if ( USE_REG ) begin : ff_1764
        reg   lut_1764_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1764_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1764_ff <= lut_1764_out;
            end
        end
        
        assign out_data[1764] = lut_1764_ff;
    end
    else begin : no_ff_1764
        assign out_data[1764] = lut_1764_out;
    end
    endgenerate
    
    
    
    // LUT : 1765
    wire [63:0] lut_1765_table = 64'b1111111111011100110111111101110011111111110111001101111111011100;
    wire [5:0] lut_1765_select = {
                             in_data[770],
                             in_data[617],
                             in_data[717],
                             in_data[178],
                             in_data[716],
                             in_data[96]};
    
    wire lut_1765_out = lut_1765_table[lut_1765_select];
    
    generate
    if ( USE_REG ) begin : ff_1765
        reg   lut_1765_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1765_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1765_ff <= lut_1765_out;
            end
        end
        
        assign out_data[1765] = lut_1765_ff;
    end
    else begin : no_ff_1765
        assign out_data[1765] = lut_1765_out;
    end
    endgenerate
    
    
    
    // LUT : 1766
    wire [63:0] lut_1766_table = 64'b0100000001000000010000000000000011010101110101011101010111010101;
    wire [5:0] lut_1766_select = {
                             in_data[709],
                             in_data[780],
                             in_data[89],
                             in_data[478],
                             in_data[13],
                             in_data[284]};
    
    wire lut_1766_out = lut_1766_table[lut_1766_select];
    
    generate
    if ( USE_REG ) begin : ff_1766
        reg   lut_1766_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1766_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1766_ff <= lut_1766_out;
            end
        end
        
        assign out_data[1766] = lut_1766_ff;
    end
    else begin : no_ff_1766
        assign out_data[1766] = lut_1766_out;
    end
    endgenerate
    
    
    
    // LUT : 1767
    wire [63:0] lut_1767_table = 64'b0000000000000000000000000000000010101111111111111011111111111111;
    wire [5:0] lut_1767_select = {
                             in_data[379],
                             in_data[419],
                             in_data[141],
                             in_data[90],
                             in_data[450],
                             in_data[655]};
    
    wire lut_1767_out = lut_1767_table[lut_1767_select];
    
    generate
    if ( USE_REG ) begin : ff_1767
        reg   lut_1767_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1767_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1767_ff <= lut_1767_out;
            end
        end
        
        assign out_data[1767] = lut_1767_ff;
    end
    else begin : no_ff_1767
        assign out_data[1767] = lut_1767_out;
    end
    endgenerate
    
    
    
    // LUT : 1768
    wire [63:0] lut_1768_table = 64'b1110111011101110111011101110111011111110111111101111111011111110;
    wire [5:0] lut_1768_select = {
                             in_data[65],
                             in_data[80],
                             in_data[589],
                             in_data[466],
                             in_data[341],
                             in_data[101]};
    
    wire lut_1768_out = lut_1768_table[lut_1768_select];
    
    generate
    if ( USE_REG ) begin : ff_1768
        reg   lut_1768_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1768_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1768_ff <= lut_1768_out;
            end
        end
        
        assign out_data[1768] = lut_1768_ff;
    end
    else begin : no_ff_1768
        assign out_data[1768] = lut_1768_out;
    end
    endgenerate
    
    
    
    // LUT : 1769
    wire [63:0] lut_1769_table = 64'b1111111100000000111111110000000011111111000000001111111110000000;
    wire [5:0] lut_1769_select = {
                             in_data[470],
                             in_data[234],
                             in_data[545],
                             in_data[534],
                             in_data[56],
                             in_data[552]};
    
    wire lut_1769_out = lut_1769_table[lut_1769_select];
    
    generate
    if ( USE_REG ) begin : ff_1769
        reg   lut_1769_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1769_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1769_ff <= lut_1769_out;
            end
        end
        
        assign out_data[1769] = lut_1769_ff;
    end
    else begin : no_ff_1769
        assign out_data[1769] = lut_1769_out;
    end
    endgenerate
    
    
    
    // LUT : 1770
    wire [63:0] lut_1770_table = 64'b0000000000000000000000000000000000000100000001000111111101111111;
    wire [5:0] lut_1770_select = {
                             in_data[628],
                             in_data[72],
                             in_data[646],
                             in_data[387],
                             in_data[373],
                             in_data[431]};
    
    wire lut_1770_out = lut_1770_table[lut_1770_select];
    
    generate
    if ( USE_REG ) begin : ff_1770
        reg   lut_1770_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1770_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1770_ff <= lut_1770_out;
            end
        end
        
        assign out_data[1770] = lut_1770_ff;
    end
    else begin : no_ff_1770
        assign out_data[1770] = lut_1770_out;
    end
    endgenerate
    
    
    
    // LUT : 1771
    wire [63:0] lut_1771_table = 64'b1111111111110000111111110000000011111111111100001111111111100000;
    wire [5:0] lut_1771_select = {
                             in_data[619],
                             in_data[39],
                             in_data[436],
                             in_data[496],
                             in_data[83],
                             in_data[169]};
    
    wire lut_1771_out = lut_1771_table[lut_1771_select];
    
    generate
    if ( USE_REG ) begin : ff_1771
        reg   lut_1771_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1771_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1771_ff <= lut_1771_out;
            end
        end
        
        assign out_data[1771] = lut_1771_ff;
    end
    else begin : no_ff_1771
        assign out_data[1771] = lut_1771_out;
    end
    endgenerate
    
    
    
    // LUT : 1772
    wire [63:0] lut_1772_table = 64'b0000000010101010101010101010101000000000101010001010101010101010;
    wire [5:0] lut_1772_select = {
                             in_data[280],
                             in_data[663],
                             in_data[651],
                             in_data[200],
                             in_data[760],
                             in_data[385]};
    
    wire lut_1772_out = lut_1772_table[lut_1772_select];
    
    generate
    if ( USE_REG ) begin : ff_1772
        reg   lut_1772_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1772_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1772_ff <= lut_1772_out;
            end
        end
        
        assign out_data[1772] = lut_1772_ff;
    end
    else begin : no_ff_1772
        assign out_data[1772] = lut_1772_out;
    end
    endgenerate
    
    
    
    // LUT : 1773
    wire [63:0] lut_1773_table = 64'b1100110011000000111111001110100011001100110000001111110011111000;
    wire [5:0] lut_1773_select = {
                             in_data[17],
                             in_data[276],
                             in_data[218],
                             in_data[272],
                             in_data[159],
                             in_data[253]};
    
    wire lut_1773_out = lut_1773_table[lut_1773_select];
    
    generate
    if ( USE_REG ) begin : ff_1773
        reg   lut_1773_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1773_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1773_ff <= lut_1773_out;
            end
        end
        
        assign out_data[1773] = lut_1773_ff;
    end
    else begin : no_ff_1773
        assign out_data[1773] = lut_1773_out;
    end
    endgenerate
    
    
    
    // LUT : 1774
    wire [63:0] lut_1774_table = 64'b1111111111001100111111111000110011111111000010001111111100001000;
    wire [5:0] lut_1774_select = {
                             in_data[523],
                             in_data[279],
                             in_data[412],
                             in_data[165],
                             in_data[486],
                             in_data[746]};
    
    wire lut_1774_out = lut_1774_table[lut_1774_select];
    
    generate
    if ( USE_REG ) begin : ff_1774
        reg   lut_1774_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1774_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1774_ff <= lut_1774_out;
            end
        end
        
        assign out_data[1774] = lut_1774_ff;
    end
    else begin : no_ff_1774
        assign out_data[1774] = lut_1774_out;
    end
    endgenerate
    
    
    
    // LUT : 1775
    wire [63:0] lut_1775_table = 64'b0000000001000100000000000100010001000101110111010100010011011101;
    wire [5:0] lut_1775_select = {
                             in_data[206],
                             in_data[20],
                             in_data[255],
                             in_data[335],
                             in_data[692],
                             in_data[521]};
    
    wire lut_1775_out = lut_1775_table[lut_1775_select];
    
    generate
    if ( USE_REG ) begin : ff_1775
        reg   lut_1775_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1775_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1775_ff <= lut_1775_out;
            end
        end
        
        assign out_data[1775] = lut_1775_ff;
    end
    else begin : no_ff_1775
        assign out_data[1775] = lut_1775_out;
    end
    endgenerate
    
    
    
    // LUT : 1776
    wire [63:0] lut_1776_table = 64'b1111001111110011111100111111111110110000101100001111000011110000;
    wire [5:0] lut_1776_select = {
                             in_data[681],
                             in_data[113],
                             in_data[0],
                             in_data[596],
                             in_data[591],
                             in_data[47]};
    
    wire lut_1776_out = lut_1776_table[lut_1776_select];
    
    generate
    if ( USE_REG ) begin : ff_1776
        reg   lut_1776_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1776_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1776_ff <= lut_1776_out;
            end
        end
        
        assign out_data[1776] = lut_1776_ff;
    end
    else begin : no_ff_1776
        assign out_data[1776] = lut_1776_out;
    end
    endgenerate
    
    
    
    // LUT : 1777
    wire [63:0] lut_1777_table = 64'b1111111111111111000011110000111111111111111111110000000000001000;
    wire [5:0] lut_1777_select = {
                             in_data[508],
                             in_data[127],
                             in_data[448],
                             in_data[177],
                             in_data[82],
                             in_data[64]};
    
    wire lut_1777_out = lut_1777_table[lut_1777_select];
    
    generate
    if ( USE_REG ) begin : ff_1777
        reg   lut_1777_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1777_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1777_ff <= lut_1777_out;
            end
        end
        
        assign out_data[1777] = lut_1777_ff;
    end
    else begin : no_ff_1777
        assign out_data[1777] = lut_1777_out;
    end
    endgenerate
    
    
    
    // LUT : 1778
    wire [63:0] lut_1778_table = 64'b1100110000000000111111111100110011111111110011001111111111111101;
    wire [5:0] lut_1778_select = {
                             in_data[635],
                             in_data[776],
                             in_data[365],
                             in_data[22],
                             in_data[145],
                             in_data[752]};
    
    wire lut_1778_out = lut_1778_table[lut_1778_select];
    
    generate
    if ( USE_REG ) begin : ff_1778
        reg   lut_1778_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1778_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1778_ff <= lut_1778_out;
            end
        end
        
        assign out_data[1778] = lut_1778_ff;
    end
    else begin : no_ff_1778
        assign out_data[1778] = lut_1778_out;
    end
    endgenerate
    
    
    
    // LUT : 1779
    wire [63:0] lut_1779_table = 64'b1010101010101010111111111111111110101010101010101111111111111111;
    wire [5:0] lut_1779_select = {
                             in_data[761],
                             in_data[342],
                             in_data[35],
                             in_data[140],
                             in_data[362],
                             in_data[395]};
    
    wire lut_1779_out = lut_1779_table[lut_1779_select];
    
    generate
    if ( USE_REG ) begin : ff_1779
        reg   lut_1779_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1779_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1779_ff <= lut_1779_out;
            end
        end
        
        assign out_data[1779] = lut_1779_ff;
    end
    else begin : no_ff_1779
        assign out_data[1779] = lut_1779_out;
    end
    endgenerate
    
    
    
    // LUT : 1780
    wire [63:0] lut_1780_table = 64'b1111110011111100111110001111100011110000111100001111000011110000;
    wire [5:0] lut_1780_select = {
                             in_data[433],
                             in_data[722],
                             in_data[281],
                             in_data[490],
                             in_data[77],
                             in_data[727]};
    
    wire lut_1780_out = lut_1780_table[lut_1780_select];
    
    generate
    if ( USE_REG ) begin : ff_1780
        reg   lut_1780_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1780_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1780_ff <= lut_1780_out;
            end
        end
        
        assign out_data[1780] = lut_1780_ff;
    end
    else begin : no_ff_1780
        assign out_data[1780] = lut_1780_out;
    end
    endgenerate
    
    
    
    // LUT : 1781
    wire [63:0] lut_1781_table = 64'b0000000011001100000000001111110000010000110111000001000011111101;
    wire [5:0] lut_1781_select = {
                             in_data[299],
                             in_data[346],
                             in_data[156],
                             in_data[745],
                             in_data[410],
                             in_data[453]};
    
    wire lut_1781_out = lut_1781_table[lut_1781_select];
    
    generate
    if ( USE_REG ) begin : ff_1781
        reg   lut_1781_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1781_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1781_ff <= lut_1781_out;
            end
        end
        
        assign out_data[1781] = lut_1781_ff;
    end
    else begin : no_ff_1781
        assign out_data[1781] = lut_1781_out;
    end
    endgenerate
    
    
    
    // LUT : 1782
    wire [63:0] lut_1782_table = 64'b1111111111111111101010101010101011111111111111111010101010101010;
    wire [5:0] lut_1782_select = {
                             in_data[654],
                             in_data[277],
                             in_data[616],
                             in_data[701],
                             in_data[476],
                             in_data[404]};
    
    wire lut_1782_out = lut_1782_table[lut_1782_select];
    
    generate
    if ( USE_REG ) begin : ff_1782
        reg   lut_1782_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1782_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1782_ff <= lut_1782_out;
            end
        end
        
        assign out_data[1782] = lut_1782_ff;
    end
    else begin : no_ff_1782
        assign out_data[1782] = lut_1782_out;
    end
    endgenerate
    
    
    
    // LUT : 1783
    wire [63:0] lut_1783_table = 64'b1111011111111111000001010000010101010111111101110000010100000101;
    wire [5:0] lut_1783_select = {
                             in_data[586],
                             in_data[537],
                             in_data[759],
                             in_data[216],
                             in_data[336],
                             in_data[339]};
    
    wire lut_1783_out = lut_1783_table[lut_1783_select];
    
    generate
    if ( USE_REG ) begin : ff_1783
        reg   lut_1783_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1783_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1783_ff <= lut_1783_out;
            end
        end
        
        assign out_data[1783] = lut_1783_ff;
    end
    else begin : no_ff_1783
        assign out_data[1783] = lut_1783_out;
    end
    endgenerate
    
    
    
    // LUT : 1784
    wire [63:0] lut_1784_table = 64'b0000000000000000000000000000010100000000000001010000000000010101;
    wire [5:0] lut_1784_select = {
                             in_data[653],
                             in_data[71],
                             in_data[501],
                             in_data[312],
                             in_data[16],
                             in_data[126]};
    
    wire lut_1784_out = lut_1784_table[lut_1784_select];
    
    generate
    if ( USE_REG ) begin : ff_1784
        reg   lut_1784_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1784_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1784_ff <= lut_1784_out;
            end
        end
        
        assign out_data[1784] = lut_1784_ff;
    end
    else begin : no_ff_1784
        assign out_data[1784] = lut_1784_out;
    end
    endgenerate
    
    
    
    // LUT : 1785
    wire [63:0] lut_1785_table = 64'b1111111010101010101011101010101011111101110010001111110111001000;
    wire [5:0] lut_1785_select = {
                             in_data[353],
                             in_data[548],
                             in_data[454],
                             in_data[622],
                             in_data[355],
                             in_data[377]};
    
    wire lut_1785_out = lut_1785_table[lut_1785_select];
    
    generate
    if ( USE_REG ) begin : ff_1785
        reg   lut_1785_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1785_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1785_ff <= lut_1785_out;
            end
        end
        
        assign out_data[1785] = lut_1785_ff;
    end
    else begin : no_ff_1785
        assign out_data[1785] = lut_1785_out;
    end
    endgenerate
    
    
    
    // LUT : 1786
    wire [63:0] lut_1786_table = 64'b1111111111111111111100001111000011111111111111111111000011110000;
    wire [5:0] lut_1786_select = {
                             in_data[706],
                             in_data[693],
                             in_data[477],
                             in_data[427],
                             in_data[451],
                             in_data[543]};
    
    wire lut_1786_out = lut_1786_table[lut_1786_select];
    
    generate
    if ( USE_REG ) begin : ff_1786
        reg   lut_1786_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1786_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1786_ff <= lut_1786_out;
            end
        end
        
        assign out_data[1786] = lut_1786_ff;
    end
    else begin : no_ff_1786
        assign out_data[1786] = lut_1786_out;
    end
    endgenerate
    
    
    
    // LUT : 1787
    wire [63:0] lut_1787_table = 64'b0001000100010001000100010001000100000000000000000000000000000000;
    wire [5:0] lut_1787_select = {
                             in_data[509],
                             in_data[779],
                             in_data[615],
                             in_data[732],
                             in_data[713],
                             in_data[720]};
    
    wire lut_1787_out = lut_1787_table[lut_1787_select];
    
    generate
    if ( USE_REG ) begin : ff_1787
        reg   lut_1787_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1787_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1787_ff <= lut_1787_out;
            end
        end
        
        assign out_data[1787] = lut_1787_ff;
    end
    else begin : no_ff_1787
        assign out_data[1787] = lut_1787_out;
    end
    endgenerate
    
    
    
    // LUT : 1788
    wire [63:0] lut_1788_table = 64'b0101111101011111000000110000000101010101010101010000010000000100;
    wire [5:0] lut_1788_select = {
                             in_data[597],
                             in_data[291],
                             in_data[43],
                             in_data[129],
                             in_data[155],
                             in_data[210]};
    
    wire lut_1788_out = lut_1788_table[lut_1788_select];
    
    generate
    if ( USE_REG ) begin : ff_1788
        reg   lut_1788_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1788_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1788_ff <= lut_1788_out;
            end
        end
        
        assign out_data[1788] = lut_1788_ff;
    end
    else begin : no_ff_1788
        assign out_data[1788] = lut_1788_out;
    end
    endgenerate
    
    
    
    // LUT : 1789
    wire [63:0] lut_1789_table = 64'b0000000010100000000011111111111100000000101000100000111111111111;
    wire [5:0] lut_1789_select = {
                             in_data[718],
                             in_data[462],
                             in_data[603],
                             in_data[624],
                             in_data[421],
                             in_data[269]};
    
    wire lut_1789_out = lut_1789_table[lut_1789_select];
    
    generate
    if ( USE_REG ) begin : ff_1789
        reg   lut_1789_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1789_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1789_ff <= lut_1789_out;
            end
        end
        
        assign out_data[1789] = lut_1789_ff;
    end
    else begin : no_ff_1789
        assign out_data[1789] = lut_1789_out;
    end
    endgenerate
    
    
    
    // LUT : 1790
    wire [63:0] lut_1790_table = 64'b0000111100001110000011110000111001011111000011000101111101001100;
    wire [5:0] lut_1790_select = {
                             in_data[181],
                             in_data[700],
                             in_data[636],
                             in_data[292],
                             in_data[459],
                             in_data[122]};
    
    wire lut_1790_out = lut_1790_table[lut_1790_select];
    
    generate
    if ( USE_REG ) begin : ff_1790
        reg   lut_1790_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1790_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1790_ff <= lut_1790_out;
            end
        end
        
        assign out_data[1790] = lut_1790_ff;
    end
    else begin : no_ff_1790
        assign out_data[1790] = lut_1790_out;
    end
    endgenerate
    
    
    
    // LUT : 1791
    wire [63:0] lut_1791_table = 64'b1100111111111111110011111111111100001111010011110000111111001111;
    wire [5:0] lut_1791_select = {
                             in_data[707],
                             in_data[782],
                             in_data[660],
                             in_data[544],
                             in_data[743],
                             in_data[224]};
    
    wire lut_1791_out = lut_1791_table[lut_1791_select];
    
    generate
    if ( USE_REG ) begin : ff_1791
        reg   lut_1791_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1791_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1791_ff <= lut_1791_out;
            end
        end
        
        assign out_data[1791] = lut_1791_ff;
    end
    else begin : no_ff_1791
        assign out_data[1791] = lut_1791_out;
    end
    endgenerate
    
    
    
    // LUT : 1792
    wire [63:0] lut_1792_table = 64'b1111111111011101111111111101110011111111110111011111111111001100;
    wire [5:0] lut_1792_select = {
                             in_data[30],
                             in_data[176],
                             in_data[358],
                             in_data[41],
                             in_data[97],
                             in_data[323]};
    
    wire lut_1792_out = lut_1792_table[lut_1792_select];
    
    generate
    if ( USE_REG ) begin : ff_1792
        reg   lut_1792_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1792_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1792_ff <= lut_1792_out;
            end
        end
        
        assign out_data[1792] = lut_1792_ff;
    end
    else begin : no_ff_1792
        assign out_data[1792] = lut_1792_out;
    end
    endgenerate
    
    
    
    // LUT : 1793
    wire [63:0] lut_1793_table = 64'b1111001111111011011100111111111100110010111000000111000111111111;
    wire [5:0] lut_1793_select = {
                             in_data[131],
                             in_data[266],
                             in_data[347],
                             in_data[73],
                             in_data[300],
                             in_data[607]};
    
    wire lut_1793_out = lut_1793_table[lut_1793_select];
    
    generate
    if ( USE_REG ) begin : ff_1793
        reg   lut_1793_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1793_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1793_ff <= lut_1793_out;
            end
        end
        
        assign out_data[1793] = lut_1793_ff;
    end
    else begin : no_ff_1793
        assign out_data[1793] = lut_1793_out;
    end
    endgenerate
    
    
    
    // LUT : 1794
    wire [63:0] lut_1794_table = 64'b0000000000001111000000000000111100000000000011110000000000101111;
    wire [5:0] lut_1794_select = {
                             in_data[50],
                             in_data[143],
                             in_data[371],
                             in_data[485],
                             in_data[270],
                             in_data[256]};
    
    wire lut_1794_out = lut_1794_table[lut_1794_select];
    
    generate
    if ( USE_REG ) begin : ff_1794
        reg   lut_1794_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1794_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1794_ff <= lut_1794_out;
            end
        end
        
        assign out_data[1794] = lut_1794_ff;
    end
    else begin : no_ff_1794
        assign out_data[1794] = lut_1794_out;
    end
    endgenerate
    
    
    
    // LUT : 1795
    wire [63:0] lut_1795_table = 64'b0010111100101111001010110010101100001011000010110000101100001011;
    wire [5:0] lut_1795_select = {
                             in_data[108],
                             in_data[76],
                             in_data[364],
                             in_data[593],
                             in_data[735],
                             in_data[777]};
    
    wire lut_1795_out = lut_1795_table[lut_1795_select];
    
    generate
    if ( USE_REG ) begin : ff_1795
        reg   lut_1795_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1795_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1795_ff <= lut_1795_out;
            end
        end
        
        assign out_data[1795] = lut_1795_ff;
    end
    else begin : no_ff_1795
        assign out_data[1795] = lut_1795_out;
    end
    endgenerate
    
    
    
    // LUT : 1796
    wire [63:0] lut_1796_table = 64'b1111111110101110111011111010111011111111101010101111111110101110;
    wire [5:0] lut_1796_select = {
                             in_data[432],
                             in_data[370],
                             in_data[748],
                             in_data[133],
                             in_data[356],
                             in_data[632]};
    
    wire lut_1796_out = lut_1796_table[lut_1796_select];
    
    generate
    if ( USE_REG ) begin : ff_1796
        reg   lut_1796_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1796_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1796_ff <= lut_1796_out;
            end
        end
        
        assign out_data[1796] = lut_1796_ff;
    end
    else begin : no_ff_1796
        assign out_data[1796] = lut_1796_out;
    end
    endgenerate
    
    
    
    // LUT : 1797
    wire [63:0] lut_1797_table = 64'b0000000000000000000100010001000000010000000000010001000100010001;
    wire [5:0] lut_1797_select = {
                             in_data[480],
                             in_data[457],
                             in_data[763],
                             in_data[60],
                             in_data[400],
                             in_data[584]};
    
    wire lut_1797_out = lut_1797_table[lut_1797_select];
    
    generate
    if ( USE_REG ) begin : ff_1797
        reg   lut_1797_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1797_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1797_ff <= lut_1797_out;
            end
        end
        
        assign out_data[1797] = lut_1797_ff;
    end
    else begin : no_ff_1797
        assign out_data[1797] = lut_1797_out;
    end
    endgenerate
    
    
    
    // LUT : 1798
    wire [63:0] lut_1798_table = 64'b0000000000000000000000010000000100000000000000000000000100000001;
    wire [5:0] lut_1798_select = {
                             in_data[767],
                             in_data[705],
                             in_data[144],
                             in_data[104],
                             in_data[229],
                             in_data[188]};
    
    wire lut_1798_out = lut_1798_table[lut_1798_select];
    
    generate
    if ( USE_REG ) begin : ff_1798
        reg   lut_1798_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1798_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1798_ff <= lut_1798_out;
            end
        end
        
        assign out_data[1798] = lut_1798_ff;
    end
    else begin : no_ff_1798
        assign out_data[1798] = lut_1798_out;
    end
    endgenerate
    
    
    
    // LUT : 1799
    wire [63:0] lut_1799_table = 64'b1111111111001100111111111100110011111111111111111111111111111111;
    wire [5:0] lut_1799_select = {
                             in_data[407],
                             in_data[446],
                             in_data[106],
                             in_data[51],
                             in_data[528],
                             in_data[734]};
    
    wire lut_1799_out = lut_1799_table[lut_1799_select];
    
    generate
    if ( USE_REG ) begin : ff_1799
        reg   lut_1799_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1799_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1799_ff <= lut_1799_out;
            end
        end
        
        assign out_data[1799] = lut_1799_ff;
    end
    else begin : no_ff_1799
        assign out_data[1799] = lut_1799_out;
    end
    endgenerate
    
    
    
    // LUT : 1800
    wire [63:0] lut_1800_table = 64'b1100110111001101110011011100110101001101010011011100110111001101;
    wire [5:0] lut_1800_select = {
                             in_data[729],
                             in_data[420],
                             in_data[618],
                             in_data[295],
                             in_data[426],
                             in_data[467]};
    
    wire lut_1800_out = lut_1800_table[lut_1800_select];
    
    generate
    if ( USE_REG ) begin : ff_1800
        reg   lut_1800_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1800_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1800_ff <= lut_1800_out;
            end
        end
        
        assign out_data[1800] = lut_1800_ff;
    end
    else begin : no_ff_1800
        assign out_data[1800] = lut_1800_out;
    end
    endgenerate
    
    
    
    // LUT : 1801
    wire [63:0] lut_1801_table = 64'b1011101110101010101110111010101010111011101010101011101110101010;
    wire [5:0] lut_1801_select = {
                             in_data[728],
                             in_data[125],
                             in_data[368],
                             in_data[723],
                             in_data[105],
                             in_data[315]};
    
    wire lut_1801_out = lut_1801_table[lut_1801_select];
    
    generate
    if ( USE_REG ) begin : ff_1801
        reg   lut_1801_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1801_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1801_ff <= lut_1801_out;
            end
        end
        
        assign out_data[1801] = lut_1801_ff;
    end
    else begin : no_ff_1801
        assign out_data[1801] = lut_1801_out;
    end
    endgenerate
    
    
    
    // LUT : 1802
    wire [63:0] lut_1802_table = 64'b1100110011111111010001001111111111001100111111110100010011011101;
    wire [5:0] lut_1802_select = {
                             in_data[198],
                             in_data[472],
                             in_data[98],
                             in_data[84],
                             in_data[738],
                             in_data[639]};
    
    wire lut_1802_out = lut_1802_table[lut_1802_select];
    
    generate
    if ( USE_REG ) begin : ff_1802
        reg   lut_1802_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1802_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1802_ff <= lut_1802_out;
            end
        end
        
        assign out_data[1802] = lut_1802_ff;
    end
    else begin : no_ff_1802
        assign out_data[1802] = lut_1802_out;
    end
    endgenerate
    
    
    
    // LUT : 1803
    wire [63:0] lut_1803_table = 64'b1100110111001101110011011100110100001100000010001010111010001100;
    wire [5:0] lut_1803_select = {
                             in_data[242],
                             in_data[375],
                             in_data[254],
                             in_data[573],
                             in_data[439],
                             in_data[237]};
    
    wire lut_1803_out = lut_1803_table[lut_1803_select];
    
    generate
    if ( USE_REG ) begin : ff_1803
        reg   lut_1803_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1803_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1803_ff <= lut_1803_out;
            end
        end
        
        assign out_data[1803] = lut_1803_ff;
    end
    else begin : no_ff_1803
        assign out_data[1803] = lut_1803_out;
    end
    endgenerate
    
    
    
    // LUT : 1804
    wire [63:0] lut_1804_table = 64'b1111010111110011111111111111001111001100110011001100110011000100;
    wire [5:0] lut_1804_select = {
                             in_data[240],
                             in_data[691],
                             in_data[482],
                             in_data[334],
                             in_data[296],
                             in_data[79]};
    
    wire lut_1804_out = lut_1804_table[lut_1804_select];
    
    generate
    if ( USE_REG ) begin : ff_1804
        reg   lut_1804_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1804_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1804_ff <= lut_1804_out;
            end
        end
        
        assign out_data[1804] = lut_1804_ff;
    end
    else begin : no_ff_1804
        assign out_data[1804] = lut_1804_out;
    end
    endgenerate
    
    
    
    // LUT : 1805
    wire [63:0] lut_1805_table = 64'b1111111111111111111111111111111111101100111111101110110011111110;
    wire [5:0] lut_1805_select = {
                             in_data[100],
                             in_data[172],
                             in_data[381],
                             in_data[652],
                             in_data[468],
                             in_data[598]};
    
    wire lut_1805_out = lut_1805_table[lut_1805_select];
    
    generate
    if ( USE_REG ) begin : ff_1805
        reg   lut_1805_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1805_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1805_ff <= lut_1805_out;
            end
        end
        
        assign out_data[1805] = lut_1805_ff;
    end
    else begin : no_ff_1805
        assign out_data[1805] = lut_1805_out;
    end
    endgenerate
    
    
    
    // LUT : 1806
    wire [63:0] lut_1806_table = 64'b1111000011110000111100001111000011111111111110101111101011111010;
    wire [5:0] lut_1806_select = {
                             in_data[241],
                             in_data[63],
                             in_data[563],
                             in_data[320],
                             in_data[48],
                             in_data[415]};
    
    wire lut_1806_out = lut_1806_table[lut_1806_select];
    
    generate
    if ( USE_REG ) begin : ff_1806
        reg   lut_1806_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1806_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1806_ff <= lut_1806_out;
            end
        end
        
        assign out_data[1806] = lut_1806_ff;
    end
    else begin : no_ff_1806
        assign out_data[1806] = lut_1806_out;
    end
    endgenerate
    
    
    
    // LUT : 1807
    wire [63:0] lut_1807_table = 64'b0000000000000000000000000000000011110000111111111111000011111110;
    wire [5:0] lut_1807_select = {
                             in_data[715],
                             in_data[57],
                             in_data[199],
                             in_data[512],
                             in_data[588],
                             in_data[222]};
    
    wire lut_1807_out = lut_1807_table[lut_1807_select];
    
    generate
    if ( USE_REG ) begin : ff_1807
        reg   lut_1807_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1807_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1807_ff <= lut_1807_out;
            end
        end
        
        assign out_data[1807] = lut_1807_ff;
    end
    else begin : no_ff_1807
        assign out_data[1807] = lut_1807_out;
    end
    endgenerate
    
    
    
    // LUT : 1808
    wire [63:0] lut_1808_table = 64'b0000010100000101000001010000010100000101000000000000010000000000;
    wire [5:0] lut_1808_select = {
                             in_data[434],
                             in_data[18],
                             in_data[162],
                             in_data[719],
                             in_data[764],
                             in_data[712]};
    
    wire lut_1808_out = lut_1808_table[lut_1808_select];
    
    generate
    if ( USE_REG ) begin : ff_1808
        reg   lut_1808_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1808_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1808_ff <= lut_1808_out;
            end
        end
        
        assign out_data[1808] = lut_1808_ff;
    end
    else begin : no_ff_1808
        assign out_data[1808] = lut_1808_out;
    end
    endgenerate
    
    
    
    // LUT : 1809
    wire [63:0] lut_1809_table = 64'b1111111111111111111111111111111011111111111111111111111111111110;
    wire [5:0] lut_1809_select = {
                             in_data[753],
                             in_data[46],
                             in_data[306],
                             in_data[449],
                             in_data[231],
                             in_data[282]};
    
    wire lut_1809_out = lut_1809_table[lut_1809_select];
    
    generate
    if ( USE_REG ) begin : ff_1809
        reg   lut_1809_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1809_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1809_ff <= lut_1809_out;
            end
        end
        
        assign out_data[1809] = lut_1809_ff;
    end
    else begin : no_ff_1809
        assign out_data[1809] = lut_1809_out;
    end
    endgenerate
    
    
    
    // LUT : 1810
    wire [63:0] lut_1810_table = 64'b0000000000001010000000000000101000001010010010100000101000001010;
    wire [5:0] lut_1810_select = {
                             in_data[585],
                             in_data[673],
                             in_data[696],
                             in_data[682],
                             in_data[781],
                             in_data[569]};
    
    wire lut_1810_out = lut_1810_table[lut_1810_select];
    
    generate
    if ( USE_REG ) begin : ff_1810
        reg   lut_1810_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1810_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1810_ff <= lut_1810_out;
            end
        end
        
        assign out_data[1810] = lut_1810_ff;
    end
    else begin : no_ff_1810
        assign out_data[1810] = lut_1810_out;
    end
    endgenerate
    
    
    
    // LUT : 1811
    wire [63:0] lut_1811_table = 64'b1000000000001000111111111000111010101010101010101111111110101111;
    wire [5:0] lut_1811_select = {
                             in_data[668],
                             in_data[208],
                             in_data[317],
                             in_data[128],
                             in_data[167],
                             in_data[135]};
    
    wire lut_1811_out = lut_1811_table[lut_1811_select];
    
    generate
    if ( USE_REG ) begin : ff_1811
        reg   lut_1811_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1811_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1811_ff <= lut_1811_out;
            end
        end
        
        assign out_data[1811] = lut_1811_ff;
    end
    else begin : no_ff_1811
        assign out_data[1811] = lut_1811_out;
    end
    endgenerate
    
    
    
    // LUT : 1812
    wire [63:0] lut_1812_table = 64'b0000000000000000000000000000110000000000000000000000000000000011;
    wire [5:0] lut_1812_select = {
                             in_data[123],
                             in_data[192],
                             in_data[189],
                             in_data[311],
                             in_data[95],
                             in_data[645]};
    
    wire lut_1812_out = lut_1812_table[lut_1812_select];
    
    generate
    if ( USE_REG ) begin : ff_1812
        reg   lut_1812_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1812_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1812_ff <= lut_1812_out;
            end
        end
        
        assign out_data[1812] = lut_1812_ff;
    end
    else begin : no_ff_1812
        assign out_data[1812] = lut_1812_out;
    end
    endgenerate
    
    
    
    // LUT : 1813
    wire [63:0] lut_1813_table = 64'b0101010100000000111111111111111101010101000000001111111111011111;
    wire [5:0] lut_1813_select = {
                             in_data[529],
                             in_data[577],
                             in_data[344],
                             in_data[675],
                             in_data[52],
                             in_data[316]};
    
    wire lut_1813_out = lut_1813_table[lut_1813_select];
    
    generate
    if ( USE_REG ) begin : ff_1813
        reg   lut_1813_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1813_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1813_ff <= lut_1813_out;
            end
        end
        
        assign out_data[1813] = lut_1813_ff;
    end
    else begin : no_ff_1813
        assign out_data[1813] = lut_1813_out;
    end
    endgenerate
    
    
    
    // LUT : 1814
    wire [63:0] lut_1814_table = 64'b0001011100000000000101110000000100010101000000000001010100000000;
    wire [5:0] lut_1814_select = {
                             in_data[174],
                             in_data[115],
                             in_data[498],
                             in_data[163],
                             in_data[243],
                             in_data[396]};
    
    wire lut_1814_out = lut_1814_table[lut_1814_select];
    
    generate
    if ( USE_REG ) begin : ff_1814
        reg   lut_1814_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1814_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1814_ff <= lut_1814_out;
            end
        end
        
        assign out_data[1814] = lut_1814_ff;
    end
    else begin : no_ff_1814
        assign out_data[1814] = lut_1814_out;
    end
    endgenerate
    
    
    
    // LUT : 1815
    wire [63:0] lut_1815_table = 64'b1111111111111111111111111111111100100011000000110010001100000010;
    wire [5:0] lut_1815_select = {
                             in_data[405],
                             in_data[308],
                             in_data[119],
                             in_data[630],
                             in_data[271],
                             in_data[443]};
    
    wire lut_1815_out = lut_1815_table[lut_1815_select];
    
    generate
    if ( USE_REG ) begin : ff_1815
        reg   lut_1815_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1815_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1815_ff <= lut_1815_out;
            end
        end
        
        assign out_data[1815] = lut_1815_ff;
    end
    else begin : no_ff_1815
        assign out_data[1815] = lut_1815_out;
    end
    endgenerate
    
    
    
    // LUT : 1816
    wire [63:0] lut_1816_table = 64'b0010000000110000001100001011001000110000001100101111001011111111;
    wire [5:0] lut_1816_select = {
                             in_data[416],
                             in_data[425],
                             in_data[367],
                             in_data[740],
                             in_data[553],
                             in_data[220]};
    
    wire lut_1816_out = lut_1816_table[lut_1816_select];
    
    generate
    if ( USE_REG ) begin : ff_1816
        reg   lut_1816_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1816_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1816_ff <= lut_1816_out;
            end
        end
        
        assign out_data[1816] = lut_1816_ff;
    end
    else begin : no_ff_1816
        assign out_data[1816] = lut_1816_out;
    end
    endgenerate
    
    
    
    // LUT : 1817
    wire [63:0] lut_1817_table = 64'b0000111100001111111111111111001001111111000111111111000000110000;
    wire [5:0] lut_1817_select = {
                             in_data[575],
                             in_data[578],
                             in_data[749],
                             in_data[235],
                             in_data[305],
                             in_data[139]};
    
    wire lut_1817_out = lut_1817_table[lut_1817_select];
    
    generate
    if ( USE_REG ) begin : ff_1817
        reg   lut_1817_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1817_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1817_ff <= lut_1817_out;
            end
        end
        
        assign out_data[1817] = lut_1817_ff;
    end
    else begin : no_ff_1817
        assign out_data[1817] = lut_1817_out;
    end
    endgenerate
    
    
    
    // LUT : 1818
    wire [63:0] lut_1818_table = 64'b1111111100001111111111110000000011111111000011110111111100000000;
    wire [5:0] lut_1818_select = {
                             in_data[58],
                             in_data[680],
                             in_data[481],
                             in_data[313],
                             in_data[765],
                             in_data[168]};
    
    wire lut_1818_out = lut_1818_table[lut_1818_select];
    
    generate
    if ( USE_REG ) begin : ff_1818
        reg   lut_1818_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1818_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1818_ff <= lut_1818_out;
            end
        end
        
        assign out_data[1818] = lut_1818_ff;
    end
    else begin : no_ff_1818
        assign out_data[1818] = lut_1818_out;
    end
    endgenerate
    
    
    
    // LUT : 1819
    wire [63:0] lut_1819_table = 64'b0000000000000000000010100000000001010000010111110101000101011111;
    wire [5:0] lut_1819_select = {
                             in_data[319],
                             in_data[34],
                             in_data[99],
                             in_data[348],
                             in_data[783],
                             in_data[160]};
    
    wire lut_1819_out = lut_1819_table[lut_1819_select];
    
    generate
    if ( USE_REG ) begin : ff_1819
        reg   lut_1819_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1819_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1819_ff <= lut_1819_out;
            end
        end
        
        assign out_data[1819] = lut_1819_ff;
    end
    else begin : no_ff_1819
        assign out_data[1819] = lut_1819_out;
    end
    endgenerate
    
    
    
    // LUT : 1820
    wire [63:0] lut_1820_table = 64'b1011111100001111101011110000111100101111000011110010111100001010;
    wire [5:0] lut_1820_select = {
                             in_data[211],
                             in_data[646],
                             in_data[741],
                             in_data[686],
                             in_data[32],
                             in_data[650]};
    
    wire lut_1820_out = lut_1820_table[lut_1820_select];
    
    generate
    if ( USE_REG ) begin : ff_1820
        reg   lut_1820_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1820_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1820_ff <= lut_1820_out;
            end
        end
        
        assign out_data[1820] = lut_1820_ff;
    end
    else begin : no_ff_1820
        assign out_data[1820] = lut_1820_out;
    end
    endgenerate
    
    
    
    // LUT : 1821
    wire [63:0] lut_1821_table = 64'b0000110001001100010011000000110011001111110011111100111111001100;
    wire [5:0] lut_1821_select = {
                             in_data[738],
                             in_data[360],
                             in_data[497],
                             in_data[739],
                             in_data[97],
                             in_data[337]};
    
    wire lut_1821_out = lut_1821_table[lut_1821_select];
    
    generate
    if ( USE_REG ) begin : ff_1821
        reg   lut_1821_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1821_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1821_ff <= lut_1821_out;
            end
        end
        
        assign out_data[1821] = lut_1821_ff;
    end
    else begin : no_ff_1821
        assign out_data[1821] = lut_1821_out;
    end
    endgenerate
    
    
    
    // LUT : 1822
    wire [63:0] lut_1822_table = 64'b1111110011111111111111001111111100000000111100000000000011110000;
    wire [5:0] lut_1822_select = {
                             in_data[464],
                             in_data[281],
                             in_data[297],
                             in_data[133],
                             in_data[435],
                             in_data[338]};
    
    wire lut_1822_out = lut_1822_table[lut_1822_select];
    
    generate
    if ( USE_REG ) begin : ff_1822
        reg   lut_1822_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1822_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1822_ff <= lut_1822_out;
            end
        end
        
        assign out_data[1822] = lut_1822_ff;
    end
    else begin : no_ff_1822
        assign out_data[1822] = lut_1822_out;
    end
    endgenerate
    
    
    
    // LUT : 1823
    wire [63:0] lut_1823_table = 64'b0000000000000000000000000000000011111100000000001111111101010011;
    wire [5:0] lut_1823_select = {
                             in_data[608],
                             in_data[77],
                             in_data[272],
                             in_data[342],
                             in_data[601],
                             in_data[422]};
    
    wire lut_1823_out = lut_1823_table[lut_1823_select];
    
    generate
    if ( USE_REG ) begin : ff_1823
        reg   lut_1823_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1823_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1823_ff <= lut_1823_out;
            end
        end
        
        assign out_data[1823] = lut_1823_ff;
    end
    else begin : no_ff_1823
        assign out_data[1823] = lut_1823_out;
    end
    endgenerate
    
    
    
    // LUT : 1824
    wire [63:0] lut_1824_table = 64'b1010101010101010101010101010101010101010101010101010101010100010;
    wire [5:0] lut_1824_select = {
                             in_data[286],
                             in_data[756],
                             in_data[645],
                             in_data[197],
                             in_data[190],
                             in_data[577]};
    
    wire lut_1824_out = lut_1824_table[lut_1824_select];
    
    generate
    if ( USE_REG ) begin : ff_1824
        reg   lut_1824_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1824_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1824_ff <= lut_1824_out;
            end
        end
        
        assign out_data[1824] = lut_1824_ff;
    end
    else begin : no_ff_1824
        assign out_data[1824] = lut_1824_out;
    end
    endgenerate
    
    
    
    // LUT : 1825
    wire [63:0] lut_1825_table = 64'b0101111100000000000011110000000111111111000000000000111100000101;
    wire [5:0] lut_1825_select = {
                             in_data[766],
                             in_data[481],
                             in_data[664],
                             in_data[255],
                             in_data[562],
                             in_data[269]};
    
    wire lut_1825_out = lut_1825_table[lut_1825_select];
    
    generate
    if ( USE_REG ) begin : ff_1825
        reg   lut_1825_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1825_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1825_ff <= lut_1825_out;
            end
        end
        
        assign out_data[1825] = lut_1825_ff;
    end
    else begin : no_ff_1825
        assign out_data[1825] = lut_1825_out;
    end
    endgenerate
    
    
    
    // LUT : 1826
    wire [63:0] lut_1826_table = 64'b0011000011111111111100001111111100110000111111110011000011111111;
    wire [5:0] lut_1826_select = {
                             in_data[122],
                             in_data[148],
                             in_data[428],
                             in_data[593],
                             in_data[351],
                             in_data[6]};
    
    wire lut_1826_out = lut_1826_table[lut_1826_select];
    
    generate
    if ( USE_REG ) begin : ff_1826
        reg   lut_1826_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1826_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1826_ff <= lut_1826_out;
            end
        end
        
        assign out_data[1826] = lut_1826_ff;
    end
    else begin : no_ff_1826
        assign out_data[1826] = lut_1826_out;
    end
    endgenerate
    
    
    
    // LUT : 1827
    wire [63:0] lut_1827_table = 64'b1010000000100000101110111011101110100000101000001011101110111011;
    wire [5:0] lut_1827_select = {
                             in_data[251],
                             in_data[604],
                             in_data[727],
                             in_data[401],
                             in_data[154],
                             in_data[273]};
    
    wire lut_1827_out = lut_1827_table[lut_1827_select];
    
    generate
    if ( USE_REG ) begin : ff_1827
        reg   lut_1827_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1827_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1827_ff <= lut_1827_out;
            end
        end
        
        assign out_data[1827] = lut_1827_ff;
    end
    else begin : no_ff_1827
        assign out_data[1827] = lut_1827_out;
    end
    endgenerate
    
    
    
    // LUT : 1828
    wire [63:0] lut_1828_table = 64'b1111000111110001111100011111000101010000011100000001000000010000;
    wire [5:0] lut_1828_select = {
                             in_data[632],
                             in_data[693],
                             in_data[506],
                             in_data[285],
                             in_data[93],
                             in_data[129]};
    
    wire lut_1828_out = lut_1828_table[lut_1828_select];
    
    generate
    if ( USE_REG ) begin : ff_1828
        reg   lut_1828_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1828_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1828_ff <= lut_1828_out;
            end
        end
        
        assign out_data[1828] = lut_1828_ff;
    end
    else begin : no_ff_1828
        assign out_data[1828] = lut_1828_out;
    end
    endgenerate
    
    
    
    // LUT : 1829
    wire [63:0] lut_1829_table = 64'b1111000011111111111111111111111100000000000000001110000000000000;
    wire [5:0] lut_1829_select = {
                             in_data[434],
                             in_data[314],
                             in_data[639],
                             in_data[514],
                             in_data[736],
                             in_data[50]};
    
    wire lut_1829_out = lut_1829_table[lut_1829_select];
    
    generate
    if ( USE_REG ) begin : ff_1829
        reg   lut_1829_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1829_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1829_ff <= lut_1829_out;
            end
        end
        
        assign out_data[1829] = lut_1829_ff;
    end
    else begin : no_ff_1829
        assign out_data[1829] = lut_1829_out;
    end
    endgenerate
    
    
    
    // LUT : 1830
    wire [63:0] lut_1830_table = 64'b1111111111111111111111111111111111111111111111111010001000000010;
    wire [5:0] lut_1830_select = {
                             in_data[745],
                             in_data[511],
                             in_data[700],
                             in_data[605],
                             in_data[679],
                             in_data[742]};
    
    wire lut_1830_out = lut_1830_table[lut_1830_select];
    
    generate
    if ( USE_REG ) begin : ff_1830
        reg   lut_1830_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1830_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1830_ff <= lut_1830_out;
            end
        end
        
        assign out_data[1830] = lut_1830_ff;
    end
    else begin : no_ff_1830
        assign out_data[1830] = lut_1830_out;
    end
    endgenerate
    
    
    
    // LUT : 1831
    wire [63:0] lut_1831_table = 64'b0101010101010101000100010001000001110111011101110001010100010001;
    wire [5:0] lut_1831_select = {
                             in_data[538],
                             in_data[120],
                             in_data[88],
                             in_data[28],
                             in_data[416],
                             in_data[375]};
    
    wire lut_1831_out = lut_1831_table[lut_1831_select];
    
    generate
    if ( USE_REG ) begin : ff_1831
        reg   lut_1831_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1831_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1831_ff <= lut_1831_out;
            end
        end
        
        assign out_data[1831] = lut_1831_ff;
    end
    else begin : no_ff_1831
        assign out_data[1831] = lut_1831_out;
    end
    endgenerate
    
    
    
    // LUT : 1832
    wire [63:0] lut_1832_table = 64'b0000000011111111110011101111111100000000111111110000000011111111;
    wire [5:0] lut_1832_select = {
                             in_data[218],
                             in_data[106],
                             in_data[353],
                             in_data[11],
                             in_data[669],
                             in_data[196]};
    
    wire lut_1832_out = lut_1832_table[lut_1832_select];
    
    generate
    if ( USE_REG ) begin : ff_1832
        reg   lut_1832_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1832_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1832_ff <= lut_1832_out;
            end
        end
        
        assign out_data[1832] = lut_1832_ff;
    end
    else begin : no_ff_1832
        assign out_data[1832] = lut_1832_out;
    end
    endgenerate
    
    
    
    // LUT : 1833
    wire [63:0] lut_1833_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_1833_select = {
                             in_data[673],
                             in_data[33],
                             in_data[350],
                             in_data[730],
                             in_data[665],
                             in_data[184]};
    
    wire lut_1833_out = lut_1833_table[lut_1833_select];
    
    generate
    if ( USE_REG ) begin : ff_1833
        reg   lut_1833_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1833_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1833_ff <= lut_1833_out;
            end
        end
        
        assign out_data[1833] = lut_1833_ff;
    end
    else begin : no_ff_1833
        assign out_data[1833] = lut_1833_out;
    end
    endgenerate
    
    
    
    // LUT : 1834
    wire [63:0] lut_1834_table = 64'b1111111111111111111111110111011111110111010101110111011100010001;
    wire [5:0] lut_1834_select = {
                             in_data[508],
                             in_data[535],
                             in_data[134],
                             in_data[280],
                             in_data[299],
                             in_data[261]};
    
    wire lut_1834_out = lut_1834_table[lut_1834_select];
    
    generate
    if ( USE_REG ) begin : ff_1834
        reg   lut_1834_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1834_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1834_ff <= lut_1834_out;
            end
        end
        
        assign out_data[1834] = lut_1834_ff;
    end
    else begin : no_ff_1834
        assign out_data[1834] = lut_1834_out;
    end
    endgenerate
    
    
    
    // LUT : 1835
    wire [63:0] lut_1835_table = 64'b0000000000000000000001001111111100000000000000000000000011111111;
    wire [5:0] lut_1835_select = {
                             in_data[363],
                             in_data[690],
                             in_data[748],
                             in_data[198],
                             in_data[476],
                             in_data[52]};
    
    wire lut_1835_out = lut_1835_table[lut_1835_select];
    
    generate
    if ( USE_REG ) begin : ff_1835
        reg   lut_1835_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1835_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1835_ff <= lut_1835_out;
            end
        end
        
        assign out_data[1835] = lut_1835_ff;
    end
    else begin : no_ff_1835
        assign out_data[1835] = lut_1835_out;
    end
    endgenerate
    
    
    
    // LUT : 1836
    wire [63:0] lut_1836_table = 64'b1111111111111111111110111111111111101000111111111111000011111110;
    wire [5:0] lut_1836_select = {
                             in_data[181],
                             in_data[654],
                             in_data[354],
                             in_data[99],
                             in_data[219],
                             in_data[305]};
    
    wire lut_1836_out = lut_1836_table[lut_1836_select];
    
    generate
    if ( USE_REG ) begin : ff_1836
        reg   lut_1836_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1836_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1836_ff <= lut_1836_out;
            end
        end
        
        assign out_data[1836] = lut_1836_ff;
    end
    else begin : no_ff_1836
        assign out_data[1836] = lut_1836_out;
    end
    endgenerate
    
    
    
    // LUT : 1837
    wire [63:0] lut_1837_table = 64'b0000000000000000000111110000111100000000000000000000111100001011;
    wire [5:0] lut_1837_select = {
                             in_data[277],
                             in_data[715],
                             in_data[647],
                             in_data[284],
                             in_data[763],
                             in_data[355]};
    
    wire lut_1837_out = lut_1837_table[lut_1837_select];
    
    generate
    if ( USE_REG ) begin : ff_1837
        reg   lut_1837_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1837_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1837_ff <= lut_1837_out;
            end
        end
        
        assign out_data[1837] = lut_1837_ff;
    end
    else begin : no_ff_1837
        assign out_data[1837] = lut_1837_out;
    end
    endgenerate
    
    
    
    // LUT : 1838
    wire [63:0] lut_1838_table = 64'b1101110111111101010100011101110111000100110111010000000001011101;
    wire [5:0] lut_1838_select = {
                             in_data[462],
                             in_data[150],
                             in_data[243],
                             in_data[624],
                             in_data[574],
                             in_data[372]};
    
    wire lut_1838_out = lut_1838_table[lut_1838_select];
    
    generate
    if ( USE_REG ) begin : ff_1838
        reg   lut_1838_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1838_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1838_ff <= lut_1838_out;
            end
        end
        
        assign out_data[1838] = lut_1838_ff;
    end
    else begin : no_ff_1838
        assign out_data[1838] = lut_1838_out;
    end
    endgenerate
    
    
    
    // LUT : 1839
    wire [63:0] lut_1839_table = 64'b1011101011111010111110101111101000000000111111110000000011111111;
    wire [5:0] lut_1839_select = {
                             in_data[541],
                             in_data[95],
                             in_data[318],
                             in_data[456],
                             in_data[74],
                             in_data[145]};
    
    wire lut_1839_out = lut_1839_table[lut_1839_select];
    
    generate
    if ( USE_REG ) begin : ff_1839
        reg   lut_1839_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1839_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1839_ff <= lut_1839_out;
            end
        end
        
        assign out_data[1839] = lut_1839_ff;
    end
    else begin : no_ff_1839
        assign out_data[1839] = lut_1839_out;
    end
    endgenerate
    
    
    
    // LUT : 1840
    wire [63:0] lut_1840_table = 64'b0000000000000000000000000000000000000000110011000000000011001100;
    wire [5:0] lut_1840_select = {
                             in_data[132],
                             in_data[558],
                             in_data[427],
                             in_data[10],
                             in_data[214],
                             in_data[591]};
    
    wire lut_1840_out = lut_1840_table[lut_1840_select];
    
    generate
    if ( USE_REG ) begin : ff_1840
        reg   lut_1840_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1840_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1840_ff <= lut_1840_out;
            end
        end
        
        assign out_data[1840] = lut_1840_ff;
    end
    else begin : no_ff_1840
        assign out_data[1840] = lut_1840_out;
    end
    endgenerate
    
    
    
    // LUT : 1841
    wire [63:0] lut_1841_table = 64'b0101010111101110000000000000000001010000000000001111111101000000;
    wire [5:0] lut_1841_select = {
                             in_data[439],
                             in_data[413],
                             in_data[543],
                             in_data[420],
                             in_data[747],
                             in_data[227]};
    
    wire lut_1841_out = lut_1841_table[lut_1841_select];
    
    generate
    if ( USE_REG ) begin : ff_1841
        reg   lut_1841_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1841_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1841_ff <= lut_1841_out;
            end
        end
        
        assign out_data[1841] = lut_1841_ff;
    end
    else begin : no_ff_1841
        assign out_data[1841] = lut_1841_out;
    end
    endgenerate
    
    
    
    // LUT : 1842
    wire [63:0] lut_1842_table = 64'b1111111111111111001100100010001011111111111111111011001100100000;
    wire [5:0] lut_1842_select = {
                             in_data[128],
                             in_data[271],
                             in_data[737],
                             in_data[774],
                             in_data[495],
                             in_data[705]};
    
    wire lut_1842_out = lut_1842_table[lut_1842_select];
    
    generate
    if ( USE_REG ) begin : ff_1842
        reg   lut_1842_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1842_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1842_ff <= lut_1842_out;
            end
        end
        
        assign out_data[1842] = lut_1842_ff;
    end
    else begin : no_ff_1842
        assign out_data[1842] = lut_1842_out;
    end
    endgenerate
    
    
    
    // LUT : 1843
    wire [63:0] lut_1843_table = 64'b1111010101000100111101010100010011110111010101001111111111010100;
    wire [5:0] lut_1843_select = {
                             in_data[389],
                             in_data[701],
                             in_data[220],
                             in_data[723],
                             in_data[287],
                             in_data[172]};
    
    wire lut_1843_out = lut_1843_table[lut_1843_select];
    
    generate
    if ( USE_REG ) begin : ff_1843
        reg   lut_1843_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1843_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1843_ff <= lut_1843_out;
            end
        end
        
        assign out_data[1843] = lut_1843_ff;
    end
    else begin : no_ff_1843
        assign out_data[1843] = lut_1843_out;
    end
    endgenerate
    
    
    
    // LUT : 1844
    wire [63:0] lut_1844_table = 64'b0000110000000000000011000000000001001100000000000100110000000100;
    wire [5:0] lut_1844_select = {
                             in_data[63],
                             in_data[370],
                             in_data[295],
                             in_data[620],
                             in_data[322],
                             in_data[761]};
    
    wire lut_1844_out = lut_1844_table[lut_1844_select];
    
    generate
    if ( USE_REG ) begin : ff_1844
        reg   lut_1844_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1844_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1844_ff <= lut_1844_out;
            end
        end
        
        assign out_data[1844] = lut_1844_ff;
    end
    else begin : no_ff_1844
        assign out_data[1844] = lut_1844_out;
    end
    endgenerate
    
    
    
    // LUT : 1845
    wire [63:0] lut_1845_table = 64'b0100010100000000010001010000000001010101000000000101010100000100;
    wire [5:0] lut_1845_select = {
                             in_data[300],
                             in_data[532],
                             in_data[412],
                             in_data[156],
                             in_data[388],
                             in_data[191]};
    
    wire lut_1845_out = lut_1845_table[lut_1845_select];
    
    generate
    if ( USE_REG ) begin : ff_1845
        reg   lut_1845_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1845_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1845_ff <= lut_1845_out;
            end
        end
        
        assign out_data[1845] = lut_1845_ff;
    end
    else begin : no_ff_1845
        assign out_data[1845] = lut_1845_out;
    end
    endgenerate
    
    
    
    // LUT : 1846
    wire [63:0] lut_1846_table = 64'b1100110011001100110011001100110011001100110011001101110111011100;
    wire [5:0] lut_1846_select = {
                             in_data[631],
                             in_data[451],
                             in_data[56],
                             in_data[782],
                             in_data[599],
                             in_data[253]};
    
    wire lut_1846_out = lut_1846_table[lut_1846_select];
    
    generate
    if ( USE_REG ) begin : ff_1846
        reg   lut_1846_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1846_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1846_ff <= lut_1846_out;
            end
        end
        
        assign out_data[1846] = lut_1846_ff;
    end
    else begin : no_ff_1846
        assign out_data[1846] = lut_1846_out;
    end
    endgenerate
    
    
    
    // LUT : 1847
    wire [63:0] lut_1847_table = 64'b0101010100000000010101010000000011111111000000001111111100000000;
    wire [5:0] lut_1847_select = {
                             in_data[432],
                             in_data[19],
                             in_data[468],
                             in_data[335],
                             in_data[304],
                             in_data[176]};
    
    wire lut_1847_out = lut_1847_table[lut_1847_select];
    
    generate
    if ( USE_REG ) begin : ff_1847
        reg   lut_1847_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1847_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1847_ff <= lut_1847_out;
            end
        end
        
        assign out_data[1847] = lut_1847_ff;
    end
    else begin : no_ff_1847
        assign out_data[1847] = lut_1847_out;
    end
    endgenerate
    
    
    
    // LUT : 1848
    wire [63:0] lut_1848_table = 64'b1111111100111111000011110000111100001111000011110000111100000010;
    wire [5:0] lut_1848_select = {
                             in_data[259],
                             in_data[692],
                             in_data[660],
                             in_data[596],
                             in_data[311],
                             in_data[105]};
    
    wire lut_1848_out = lut_1848_table[lut_1848_select];
    
    generate
    if ( USE_REG ) begin : ff_1848
        reg   lut_1848_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1848_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1848_ff <= lut_1848_out;
            end
        end
        
        assign out_data[1848] = lut_1848_ff;
    end
    else begin : no_ff_1848
        assign out_data[1848] = lut_1848_out;
    end
    endgenerate
    
    
    
    // LUT : 1849
    wire [63:0] lut_1849_table = 64'b1111111111111111101110111011101111111111111111110010001000100010;
    wire [5:0] lut_1849_select = {
                             in_data[173],
                             in_data[453],
                             in_data[25],
                             in_data[26],
                             in_data[662],
                             in_data[203]};
    
    wire lut_1849_out = lut_1849_table[lut_1849_select];
    
    generate
    if ( USE_REG ) begin : ff_1849
        reg   lut_1849_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1849_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1849_ff <= lut_1849_out;
            end
        end
        
        assign out_data[1849] = lut_1849_ff;
    end
    else begin : no_ff_1849
        assign out_data[1849] = lut_1849_out;
    end
    endgenerate
    
    
    
    // LUT : 1850
    wire [63:0] lut_1850_table = 64'b0100111101001111010011110100111101001101010011010100110001001100;
    wire [5:0] lut_1850_select = {
                             in_data[444],
                             in_data[523],
                             in_data[36],
                             in_data[230],
                             in_data[125],
                             in_data[248]};
    
    wire lut_1850_out = lut_1850_table[lut_1850_select];
    
    generate
    if ( USE_REG ) begin : ff_1850
        reg   lut_1850_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1850_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1850_ff <= lut_1850_out;
            end
        end
        
        assign out_data[1850] = lut_1850_ff;
    end
    else begin : no_ff_1850
        assign out_data[1850] = lut_1850_out;
    end
    endgenerate
    
    
    
    // LUT : 1851
    wire [63:0] lut_1851_table = 64'b1111111111111111001100110011001100110011001100110001000000010001;
    wire [5:0] lut_1851_select = {
                             in_data[121],
                             in_data[49],
                             in_data[15],
                             in_data[450],
                             in_data[663],
                             in_data[771]};
    
    wire lut_1851_out = lut_1851_table[lut_1851_select];
    
    generate
    if ( USE_REG ) begin : ff_1851
        reg   lut_1851_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1851_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1851_ff <= lut_1851_out;
            end
        end
        
        assign out_data[1851] = lut_1851_ff;
    end
    else begin : no_ff_1851
        assign out_data[1851] = lut_1851_out;
    end
    endgenerate
    
    
    
    // LUT : 1852
    wire [63:0] lut_1852_table = 64'b0000110011001100000011001100110000001100110011000000110001001100;
    wire [5:0] lut_1852_select = {
                             in_data[94],
                             in_data[87],
                             in_data[303],
                             in_data[595],
                             in_data[352],
                             in_data[642]};
    
    wire lut_1852_out = lut_1852_table[lut_1852_select];
    
    generate
    if ( USE_REG ) begin : ff_1852
        reg   lut_1852_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1852_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1852_ff <= lut_1852_out;
            end
        end
        
        assign out_data[1852] = lut_1852_ff;
    end
    else begin : no_ff_1852
        assign out_data[1852] = lut_1852_out;
    end
    endgenerate
    
    
    
    // LUT : 1853
    wire [63:0] lut_1853_table = 64'b0000001100110011000000000000000000111011001100110011001100110011;
    wire [5:0] lut_1853_select = {
                             in_data[429],
                             in_data[638],
                             in_data[395],
                             in_data[339],
                             in_data[136],
                             in_data[224]};
    
    wire lut_1853_out = lut_1853_table[lut_1853_select];
    
    generate
    if ( USE_REG ) begin : ff_1853
        reg   lut_1853_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1853_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1853_ff <= lut_1853_out;
            end
        end
        
        assign out_data[1853] = lut_1853_ff;
    end
    else begin : no_ff_1853
        assign out_data[1853] = lut_1853_out;
    end
    endgenerate
    
    
    
    // LUT : 1854
    wire [63:0] lut_1854_table = 64'b1111111110110011111111111011001111111111001100111111111100110011;
    wire [5:0] lut_1854_select = {
                             in_data[89],
                             in_data[589],
                             in_data[192],
                             in_data[42],
                             in_data[498],
                             in_data[91]};
    
    wire lut_1854_out = lut_1854_table[lut_1854_select];
    
    generate
    if ( USE_REG ) begin : ff_1854
        reg   lut_1854_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1854_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1854_ff <= lut_1854_out;
            end
        end
        
        assign out_data[1854] = lut_1854_ff;
    end
    else begin : no_ff_1854
        assign out_data[1854] = lut_1854_out;
    end
    endgenerate
    
    
    
    // LUT : 1855
    wire [63:0] lut_1855_table = 64'b1111111111111111111111111111111011101110111011101110111011101110;
    wire [5:0] lut_1855_select = {
                             in_data[207],
                             in_data[21],
                             in_data[617],
                             in_data[92],
                             in_data[499],
                             in_data[659]};
    
    wire lut_1855_out = lut_1855_table[lut_1855_select];
    
    generate
    if ( USE_REG ) begin : ff_1855
        reg   lut_1855_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1855_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1855_ff <= lut_1855_out;
            end
        end
        
        assign out_data[1855] = lut_1855_ff;
    end
    else begin : no_ff_1855
        assign out_data[1855] = lut_1855_out;
    end
    endgenerate
    
    
    
    // LUT : 1856
    wire [63:0] lut_1856_table = 64'b0001001100000001001100110001001100010001000000000011000100010001;
    wire [5:0] lut_1856_select = {
                             in_data[69],
                             in_data[594],
                             in_data[676],
                             in_data[661],
                             in_data[509],
                             in_data[446]};
    
    wire lut_1856_out = lut_1856_table[lut_1856_select];
    
    generate
    if ( USE_REG ) begin : ff_1856
        reg   lut_1856_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1856_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1856_ff <= lut_1856_out;
            end
        end
        
        assign out_data[1856] = lut_1856_ff;
    end
    else begin : no_ff_1856
        assign out_data[1856] = lut_1856_out;
    end
    endgenerate
    
    
    
    // LUT : 1857
    wire [63:0] lut_1857_table = 64'b1111111101010001111111110101000011111111010101011111111101010001;
    wire [5:0] lut_1857_select = {
                             in_data[38],
                             in_data[505],
                             in_data[341],
                             in_data[309],
                             in_data[306],
                             in_data[231]};
    
    wire lut_1857_out = lut_1857_table[lut_1857_select];
    
    generate
    if ( USE_REG ) begin : ff_1857
        reg   lut_1857_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1857_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1857_ff <= lut_1857_out;
            end
        end
        
        assign out_data[1857] = lut_1857_ff;
    end
    else begin : no_ff_1857
        assign out_data[1857] = lut_1857_out;
    end
    endgenerate
    
    
    
    // LUT : 1858
    wire [63:0] lut_1858_table = 64'b0001000000010000000100000011000011110111001100110011001000110011;
    wire [5:0] lut_1858_select = {
                             in_data[467],
                             in_data[379],
                             in_data[714],
                             in_data[666],
                             in_data[376],
                             in_data[159]};
    
    wire lut_1858_out = lut_1858_table[lut_1858_select];
    
    generate
    if ( USE_REG ) begin : ff_1858
        reg   lut_1858_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1858_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1858_ff <= lut_1858_out;
            end
        end
        
        assign out_data[1858] = lut_1858_ff;
    end
    else begin : no_ff_1858
        assign out_data[1858] = lut_1858_out;
    end
    endgenerate
    
    
    
    // LUT : 1859
    wire [63:0] lut_1859_table = 64'b1010101010101010101010101010101010101010101111101010101010101010;
    wire [5:0] lut_1859_select = {
                             in_data[493],
                             in_data[653],
                             in_data[502],
                             in_data[188],
                             in_data[465],
                             in_data[260]};
    
    wire lut_1859_out = lut_1859_table[lut_1859_select];
    
    generate
    if ( USE_REG ) begin : ff_1859
        reg   lut_1859_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1859_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1859_ff <= lut_1859_out;
            end
        end
        
        assign out_data[1859] = lut_1859_ff;
    end
    else begin : no_ff_1859
        assign out_data[1859] = lut_1859_out;
    end
    endgenerate
    
    
    
    // LUT : 1860
    wire [63:0] lut_1860_table = 64'b1010101010101010101010101010101010101010101010111010101000001010;
    wire [5:0] lut_1860_select = {
                             in_data[731],
                             in_data[381],
                             in_data[70],
                             in_data[152],
                             in_data[398],
                             in_data[289]};
    
    wire lut_1860_out = lut_1860_table[lut_1860_select];
    
    generate
    if ( USE_REG ) begin : ff_1860
        reg   lut_1860_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1860_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1860_ff <= lut_1860_out;
            end
        end
        
        assign out_data[1860] = lut_1860_ff;
    end
    else begin : no_ff_1860
        assign out_data[1860] = lut_1860_out;
    end
    endgenerate
    
    
    
    // LUT : 1861
    wire [63:0] lut_1861_table = 64'b1111111111111111111111111111011100000000000000000000001000000000;
    wire [5:0] lut_1861_select = {
                             in_data[328],
                             in_data[402],
                             in_data[1],
                             in_data[195],
                             in_data[107],
                             in_data[565]};
    
    wire lut_1861_out = lut_1861_table[lut_1861_select];
    
    generate
    if ( USE_REG ) begin : ff_1861
        reg   lut_1861_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1861_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1861_ff <= lut_1861_out;
            end
        end
        
        assign out_data[1861] = lut_1861_ff;
    end
    else begin : no_ff_1861
        assign out_data[1861] = lut_1861_out;
    end
    endgenerate
    
    
    
    // LUT : 1862
    wire [63:0] lut_1862_table = 64'b0000111100001011000011110000001100001111000010110000111100000011;
    wire [5:0] lut_1862_select = {
                             in_data[169],
                             in_data[115],
                             in_data[563],
                             in_data[636],
                             in_data[81],
                             in_data[171]};
    
    wire lut_1862_out = lut_1862_table[lut_1862_select];
    
    generate
    if ( USE_REG ) begin : ff_1862
        reg   lut_1862_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1862_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1862_ff <= lut_1862_out;
            end
        end
        
        assign out_data[1862] = lut_1862_ff;
    end
    else begin : no_ff_1862
        assign out_data[1862] = lut_1862_out;
    end
    endgenerate
    
    
    
    // LUT : 1863
    wire [63:0] lut_1863_table = 64'b1111111111111111111111101111110011111111111111111111111011111100;
    wire [5:0] lut_1863_select = {
                             in_data[48],
                             in_data[482],
                             in_data[540],
                             in_data[610],
                             in_data[473],
                             in_data[200]};
    
    wire lut_1863_out = lut_1863_table[lut_1863_select];
    
    generate
    if ( USE_REG ) begin : ff_1863
        reg   lut_1863_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1863_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1863_ff <= lut_1863_out;
            end
        end
        
        assign out_data[1863] = lut_1863_ff;
    end
    else begin : no_ff_1863
        assign out_data[1863] = lut_1863_out;
    end
    endgenerate
    
    
    
    // LUT : 1864
    wire [63:0] lut_1864_table = 64'b0000000000000000000000000000000000000000010101010000000000010101;
    wire [5:0] lut_1864_select = {
                             in_data[340],
                             in_data[55],
                             in_data[296],
                             in_data[770],
                             in_data[51],
                             in_data[711]};
    
    wire lut_1864_out = lut_1864_table[lut_1864_select];
    
    generate
    if ( USE_REG ) begin : ff_1864
        reg   lut_1864_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1864_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1864_ff <= lut_1864_out;
            end
        end
        
        assign out_data[1864] = lut_1864_ff;
    end
    else begin : no_ff_1864
        assign out_data[1864] = lut_1864_out;
    end
    endgenerate
    
    
    
    // LUT : 1865
    wire [63:0] lut_1865_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_1865_select = {
                             in_data[315],
                             in_data[78],
                             in_data[760],
                             in_data[123],
                             in_data[177],
                             in_data[728]};
    
    wire lut_1865_out = lut_1865_table[lut_1865_select];
    
    generate
    if ( USE_REG ) begin : ff_1865
        reg   lut_1865_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1865_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1865_ff <= lut_1865_out;
            end
        end
        
        assign out_data[1865] = lut_1865_ff;
    end
    else begin : no_ff_1865
        assign out_data[1865] = lut_1865_out;
    end
    endgenerate
    
    
    
    // LUT : 1866
    wire [63:0] lut_1866_table = 64'b0100010001000100000000000000000000010000000100010011001100010111;
    wire [5:0] lut_1866_select = {
                             in_data[626],
                             in_data[274],
                             in_data[472],
                             in_data[7],
                             in_data[635],
                             in_data[179]};
    
    wire lut_1866_out = lut_1866_table[lut_1866_select];
    
    generate
    if ( USE_REG ) begin : ff_1866
        reg   lut_1866_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1866_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1866_ff <= lut_1866_out;
            end
        end
        
        assign out_data[1866] = lut_1866_ff;
    end
    else begin : no_ff_1866
        assign out_data[1866] = lut_1866_out;
    end
    endgenerate
    
    
    
    // LUT : 1867
    wire [63:0] lut_1867_table = 64'b0000110011001101000011001100110000000000111111110000000011111110;
    wire [5:0] lut_1867_select = {
                             in_data[681],
                             in_data[588],
                             in_data[525],
                             in_data[487],
                             in_data[519],
                             in_data[699]};
    
    wire lut_1867_out = lut_1867_table[lut_1867_select];
    
    generate
    if ( USE_REG ) begin : ff_1867
        reg   lut_1867_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1867_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1867_ff <= lut_1867_out;
            end
        end
        
        assign out_data[1867] = lut_1867_ff;
    end
    else begin : no_ff_1867
        assign out_data[1867] = lut_1867_out;
    end
    endgenerate
    
    
    
    // LUT : 1868
    wire [63:0] lut_1868_table = 64'b0000101100001111000011110000111100000000000000010000010100000101;
    wire [5:0] lut_1868_select = {
                             in_data[597],
                             in_data[655],
                             in_data[552],
                             in_data[186],
                             in_data[529],
                             in_data[178]};
    
    wire lut_1868_out = lut_1868_table[lut_1868_select];
    
    generate
    if ( USE_REG ) begin : ff_1868
        reg   lut_1868_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1868_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1868_ff <= lut_1868_out;
            end
        end
        
        assign out_data[1868] = lut_1868_ff;
    end
    else begin : no_ff_1868
        assign out_data[1868] = lut_1868_out;
    end
    endgenerate
    
    
    
    // LUT : 1869
    wire [63:0] lut_1869_table = 64'b1011101110111011101100100011001110111011001110111011001100110011;
    wire [5:0] lut_1869_select = {
                             in_data[75],
                             in_data[707],
                             in_data[236],
                             in_data[232],
                             in_data[567],
                             in_data[649]};
    
    wire lut_1869_out = lut_1869_table[lut_1869_select];
    
    generate
    if ( USE_REG ) begin : ff_1869
        reg   lut_1869_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1869_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1869_ff <= lut_1869_out;
            end
        end
        
        assign out_data[1869] = lut_1869_ff;
    end
    else begin : no_ff_1869
        assign out_data[1869] = lut_1869_out;
    end
    endgenerate
    
    
    
    // LUT : 1870
    wire [63:0] lut_1870_table = 64'b0000000000000000000000000000000000000000000100010000000000010001;
    wire [5:0] lut_1870_select = {
                             in_data[202],
                             in_data[672],
                             in_data[367],
                             in_data[324],
                             in_data[722],
                             in_data[668]};
    
    wire lut_1870_out = lut_1870_table[lut_1870_select];
    
    generate
    if ( USE_REG ) begin : ff_1870
        reg   lut_1870_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1870_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1870_ff <= lut_1870_out;
            end
        end
        
        assign out_data[1870] = lut_1870_ff;
    end
    else begin : no_ff_1870
        assign out_data[1870] = lut_1870_out;
    end
    endgenerate
    
    
    
    // LUT : 1871
    wire [63:0] lut_1871_table = 64'b0000111100001111000000000000000000001111000011110000000000000100;
    wire [5:0] lut_1871_select = {
                             in_data[139],
                             in_data[718],
                             in_data[754],
                             in_data[773],
                             in_data[752],
                             in_data[22]};
    
    wire lut_1871_out = lut_1871_table[lut_1871_select];
    
    generate
    if ( USE_REG ) begin : ff_1871
        reg   lut_1871_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1871_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1871_ff <= lut_1871_out;
            end
        end
        
        assign out_data[1871] = lut_1871_ff;
    end
    else begin : no_ff_1871
        assign out_data[1871] = lut_1871_out;
    end
    endgenerate
    
    
    
    // LUT : 1872
    wire [63:0] lut_1872_table = 64'b1111101011111110111110101111111010110010111110101011001011111010;
    wire [5:0] lut_1872_select = {
                             in_data[330],
                             in_data[703],
                             in_data[262],
                             in_data[124],
                             in_data[189],
                             in_data[452]};
    
    wire lut_1872_out = lut_1872_table[lut_1872_select];
    
    generate
    if ( USE_REG ) begin : ff_1872
        reg   lut_1872_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1872_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1872_ff <= lut_1872_out;
            end
        end
        
        assign out_data[1872] = lut_1872_ff;
    end
    else begin : no_ff_1872
        assign out_data[1872] = lut_1872_out;
    end
    endgenerate
    
    
    
    // LUT : 1873
    wire [63:0] lut_1873_table = 64'b1111111110101010111111111110101011111111101010101111111110101010;
    wire [5:0] lut_1873_select = {
                             in_data[140],
                             in_data[616],
                             in_data[165],
                             in_data[16],
                             in_data[108],
                             in_data[521]};
    
    wire lut_1873_out = lut_1873_table[lut_1873_select];
    
    generate
    if ( USE_REG ) begin : ff_1873
        reg   lut_1873_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1873_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1873_ff <= lut_1873_out;
            end
        end
        
        assign out_data[1873] = lut_1873_ff;
    end
    else begin : no_ff_1873
        assign out_data[1873] = lut_1873_out;
    end
    endgenerate
    
    
    
    // LUT : 1874
    wire [63:0] lut_1874_table = 64'b0000000011111111000000001011111111111111111111110000000011111111;
    wire [5:0] lut_1874_select = {
                             in_data[440],
                             in_data[424],
                             in_data[458],
                             in_data[744],
                             in_data[533],
                             in_data[283]};
    
    wire lut_1874_out = lut_1874_table[lut_1874_select];
    
    generate
    if ( USE_REG ) begin : ff_1874
        reg   lut_1874_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1874_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1874_ff <= lut_1874_out;
            end
        end
        
        assign out_data[1874] = lut_1874_ff;
    end
    else begin : no_ff_1874
        assign out_data[1874] = lut_1874_out;
    end
    endgenerate
    
    
    
    // LUT : 1875
    wire [63:0] lut_1875_table = 64'b1111111111111111000000000101010111111111111111110000000000010000;
    wire [5:0] lut_1875_select = {
                             in_data[696],
                             in_data[378],
                             in_data[607],
                             in_data[503],
                             in_data[53],
                             in_data[347]};
    
    wire lut_1875_out = lut_1875_table[lut_1875_select];
    
    generate
    if ( USE_REG ) begin : ff_1875
        reg   lut_1875_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1875_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1875_ff <= lut_1875_out;
            end
        end
        
        assign out_data[1875] = lut_1875_ff;
    end
    else begin : no_ff_1875
        assign out_data[1875] = lut_1875_out;
    end
    endgenerate
    
    
    
    // LUT : 1876
    wire [63:0] lut_1876_table = 64'b0011000011110011000000000000000000110000111100110000000000100000;
    wire [5:0] lut_1876_select = {
                             in_data[474],
                             in_data[213],
                             in_data[709],
                             in_data[405],
                             in_data[71],
                             in_data[734]};
    
    wire lut_1876_out = lut_1876_table[lut_1876_select];
    
    generate
    if ( USE_REG ) begin : ff_1876
        reg   lut_1876_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1876_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1876_ff <= lut_1876_out;
            end
        end
        
        assign out_data[1876] = lut_1876_ff;
    end
    else begin : no_ff_1876
        assign out_data[1876] = lut_1876_out;
    end
    endgenerate
    
    
    
    // LUT : 1877
    wire [63:0] lut_1877_table = 64'b1111111111111111111111111111101111011101110111011111101111110001;
    wire [5:0] lut_1877_select = {
                             in_data[501],
                             in_data[175],
                             in_data[732],
                             in_data[500],
                             in_data[265],
                             in_data[460]};
    
    wire lut_1877_out = lut_1877_table[lut_1877_select];
    
    generate
    if ( USE_REG ) begin : ff_1877
        reg   lut_1877_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1877_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1877_ff <= lut_1877_out;
            end
        end
        
        assign out_data[1877] = lut_1877_ff;
    end
    else begin : no_ff_1877
        assign out_data[1877] = lut_1877_out;
    end
    endgenerate
    
    
    
    // LUT : 1878
    wire [63:0] lut_1878_table = 64'b0010111100001010000011110000101010101111101011110000111100001111;
    wire [5:0] lut_1878_select = {
                             in_data[72],
                             in_data[327],
                             in_data[549],
                             in_data[516],
                             in_data[222],
                             in_data[201]};
    
    wire lut_1878_out = lut_1878_table[lut_1878_select];
    
    generate
    if ( USE_REG ) begin : ff_1878
        reg   lut_1878_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1878_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1878_ff <= lut_1878_out;
            end
        end
        
        assign out_data[1878] = lut_1878_ff;
    end
    else begin : no_ff_1878
        assign out_data[1878] = lut_1878_out;
    end
    endgenerate
    
    
    
    // LUT : 1879
    wire [63:0] lut_1879_table = 64'b0000101100001010100011111000111100000010000000000000111100001111;
    wire [5:0] lut_1879_select = {
                             in_data[557],
                             in_data[247],
                             in_data[254],
                             in_data[301],
                             in_data[454],
                             in_data[582]};
    
    wire lut_1879_out = lut_1879_table[lut_1879_select];
    
    generate
    if ( USE_REG ) begin : ff_1879
        reg   lut_1879_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1879_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1879_ff <= lut_1879_out;
            end
        end
        
        assign out_data[1879] = lut_1879_ff;
    end
    else begin : no_ff_1879
        assign out_data[1879] = lut_1879_out;
    end
    endgenerate
    
    
    
    // LUT : 1880
    wire [63:0] lut_1880_table = 64'b0011000000110000101100001111000011110000111100001111000011110010;
    wire [5:0] lut_1880_select = {
                             in_data[708],
                             in_data[221],
                             in_data[380],
                             in_data[602],
                             in_data[489],
                             in_data[590]};
    
    wire lut_1880_out = lut_1880_table[lut_1880_select];
    
    generate
    if ( USE_REG ) begin : ff_1880
        reg   lut_1880_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1880_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1880_ff <= lut_1880_out;
            end
        end
        
        assign out_data[1880] = lut_1880_ff;
    end
    else begin : no_ff_1880
        assign out_data[1880] = lut_1880_out;
    end
    endgenerate
    
    
    
    // LUT : 1881
    wire [63:0] lut_1881_table = 64'b0000000000000000000000100000000011111111111011101111111101110111;
    wire [5:0] lut_1881_select = {
                             in_data[294],
                             in_data[581],
                             in_data[396],
                             in_data[54],
                             in_data[547],
                             in_data[575]};
    
    wire lut_1881_out = lut_1881_table[lut_1881_select];
    
    generate
    if ( USE_REG ) begin : ff_1881
        reg   lut_1881_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1881_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1881_ff <= lut_1881_out;
            end
        end
        
        assign out_data[1881] = lut_1881_ff;
    end
    else begin : no_ff_1881
        assign out_data[1881] = lut_1881_out;
    end
    endgenerate
    
    
    
    // LUT : 1882
    wire [63:0] lut_1882_table = 64'b0011001100000000001100110011001100110011000000000011001100110011;
    wire [5:0] lut_1882_select = {
                             in_data[674],
                             in_data[374],
                             in_data[241],
                             in_data[334],
                             in_data[470],
                             in_data[671]};
    
    wire lut_1882_out = lut_1882_table[lut_1882_select];
    
    generate
    if ( USE_REG ) begin : ff_1882
        reg   lut_1882_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1882_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1882_ff <= lut_1882_out;
            end
        end
        
        assign out_data[1882] = lut_1882_ff;
    end
    else begin : no_ff_1882
        assign out_data[1882] = lut_1882_out;
    end
    endgenerate
    
    
    
    // LUT : 1883
    wire [63:0] lut_1883_table = 64'b0000000010101011000000000010101000000000001010100000000000101010;
    wire [5:0] lut_1883_select = {
                             in_data[366],
                             in_data[757],
                             in_data[479],
                             in_data[278],
                             in_data[144],
                             in_data[657]};
    
    wire lut_1883_out = lut_1883_table[lut_1883_select];
    
    generate
    if ( USE_REG ) begin : ff_1883
        reg   lut_1883_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1883_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1883_ff <= lut_1883_out;
            end
        end
        
        assign out_data[1883] = lut_1883_ff;
    end
    else begin : no_ff_1883
        assign out_data[1883] = lut_1883_out;
    end
    endgenerate
    
    
    
    // LUT : 1884
    wire [63:0] lut_1884_table = 64'b0000000000111011000000000011111100000000111110100000000011111010;
    wire [5:0] lut_1884_select = {
                             in_data[298],
                             in_data[116],
                             in_data[471],
                             in_data[215],
                             in_data[229],
                             in_data[537]};
    
    wire lut_1884_out = lut_1884_table[lut_1884_select];
    
    generate
    if ( USE_REG ) begin : ff_1884
        reg   lut_1884_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1884_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1884_ff <= lut_1884_out;
            end
        end
        
        assign out_data[1884] = lut_1884_ff;
    end
    else begin : no_ff_1884
        assign out_data[1884] = lut_1884_out;
    end
    endgenerate
    
    
    
    // LUT : 1885
    wire [63:0] lut_1885_table = 64'b1111110011111100111111001111110000001100000011000000110000001100;
    wire [5:0] lut_1885_select = {
                             in_data[513],
                             in_data[146],
                             in_data[729],
                             in_data[386],
                             in_data[441],
                             in_data[23]};
    
    wire lut_1885_out = lut_1885_table[lut_1885_select];
    
    generate
    if ( USE_REG ) begin : ff_1885
        reg   lut_1885_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1885_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1885_ff <= lut_1885_out;
            end
        end
        
        assign out_data[1885] = lut_1885_ff;
    end
    else begin : no_ff_1885
        assign out_data[1885] = lut_1885_out;
    end
    endgenerate
    
    
    
    // LUT : 1886
    wire [63:0] lut_1886_table = 64'b1101000001010000110100010101000011010000010100001101000011010000;
    wire [5:0] lut_1886_select = {
                             in_data[759],
                             in_data[168],
                             in_data[762],
                             in_data[461],
                             in_data[687],
                             in_data[706]};
    
    wire lut_1886_out = lut_1886_table[lut_1886_select];
    
    generate
    if ( USE_REG ) begin : ff_1886
        reg   lut_1886_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1886_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1886_ff <= lut_1886_out;
            end
        end
        
        assign out_data[1886] = lut_1886_ff;
    end
    else begin : no_ff_1886
        assign out_data[1886] = lut_1886_out;
    end
    endgenerate
    
    
    
    // LUT : 1887
    wire [63:0] lut_1887_table = 64'b0000000000000000000000101000101000111011101010100011101110101110;
    wire [5:0] lut_1887_select = {
                             in_data[149],
                             in_data[187],
                             in_data[385],
                             in_data[743],
                             in_data[326],
                             in_data[358]};
    
    wire lut_1887_out = lut_1887_table[lut_1887_select];
    
    generate
    if ( USE_REG ) begin : ff_1887
        reg   lut_1887_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1887_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1887_ff <= lut_1887_out;
            end
        end
        
        assign out_data[1887] = lut_1887_ff;
    end
    else begin : no_ff_1887
        assign out_data[1887] = lut_1887_out;
    end
    endgenerate
    
    
    
    // LUT : 1888
    wire [63:0] lut_1888_table = 64'b1111111111111111000000000000000011110011111100111111111111111111;
    wire [5:0] lut_1888_select = {
                             in_data[522],
                             in_data[369],
                             in_data[447],
                             in_data[161],
                             in_data[194],
                             in_data[776]};
    
    wire lut_1888_out = lut_1888_table[lut_1888_select];
    
    generate
    if ( USE_REG ) begin : ff_1888
        reg   lut_1888_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1888_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1888_ff <= lut_1888_out;
            end
        end
        
        assign out_data[1888] = lut_1888_ff;
    end
    else begin : no_ff_1888
        assign out_data[1888] = lut_1888_out;
    end
    endgenerate
    
    
    
    // LUT : 1889
    wire [63:0] lut_1889_table = 64'b1011001110111011101110111011101110100010101000101010101010101010;
    wire [5:0] lut_1889_select = {
                             in_data[634],
                             in_data[170],
                             in_data[82],
                             in_data[554],
                             in_data[652],
                             in_data[667]};
    
    wire lut_1889_out = lut_1889_table[lut_1889_select];
    
    generate
    if ( USE_REG ) begin : ff_1889
        reg   lut_1889_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1889_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1889_ff <= lut_1889_out;
            end
        end
        
        assign out_data[1889] = lut_1889_ff;
    end
    else begin : no_ff_1889
        assign out_data[1889] = lut_1889_out;
    end
    endgenerate
    
    
    
    // LUT : 1890
    wire [63:0] lut_1890_table = 64'b0000010100001111000011110000111100000101000011110000010100001111;
    wire [5:0] lut_1890_select = {
                             in_data[46],
                             in_data[618],
                             in_data[769],
                             in_data[130],
                             in_data[308],
                             in_data[548]};
    
    wire lut_1890_out = lut_1890_table[lut_1890_select];
    
    generate
    if ( USE_REG ) begin : ff_1890
        reg   lut_1890_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1890_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1890_ff <= lut_1890_out;
            end
        end
        
        assign out_data[1890] = lut_1890_ff;
    end
    else begin : no_ff_1890
        assign out_data[1890] = lut_1890_out;
    end
    endgenerate
    
    
    
    // LUT : 1891
    wire [63:0] lut_1891_table = 64'b1010111011111111101011101111111100000000101010100000000010101010;
    wire [5:0] lut_1891_select = {
                             in_data[383],
                             in_data[58],
                             in_data[530],
                             in_data[167],
                             in_data[619],
                             in_data[67]};
    
    wire lut_1891_out = lut_1891_table[lut_1891_select];
    
    generate
    if ( USE_REG ) begin : ff_1891
        reg   lut_1891_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1891_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1891_ff <= lut_1891_out;
            end
        end
        
        assign out_data[1891] = lut_1891_ff;
    end
    else begin : no_ff_1891
        assign out_data[1891] = lut_1891_out;
    end
    endgenerate
    
    
    
    // LUT : 1892
    wire [63:0] lut_1892_table = 64'b0010111100000010001111110000001000000011000000000000001100000000;
    wire [5:0] lut_1892_select = {
                             in_data[627],
                             in_data[113],
                             in_data[320],
                             in_data[527],
                             in_data[612],
                             in_data[162]};
    
    wire lut_1892_out = lut_1892_table[lut_1892_select];
    
    generate
    if ( USE_REG ) begin : ff_1892
        reg   lut_1892_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1892_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1892_ff <= lut_1892_out;
            end
        end
        
        assign out_data[1892] = lut_1892_ff;
    end
    else begin : no_ff_1892
        assign out_data[1892] = lut_1892_out;
    end
    endgenerate
    
    
    
    // LUT : 1893
    wire [63:0] lut_1893_table = 64'b0000000000000000000111110001111100000000000000000000111100001111;
    wire [5:0] lut_1893_select = {
                             in_data[85],
                             in_data[206],
                             in_data[534],
                             in_data[406],
                             in_data[449],
                             in_data[44]};
    
    wire lut_1893_out = lut_1893_table[lut_1893_select];
    
    generate
    if ( USE_REG ) begin : ff_1893
        reg   lut_1893_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1893_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1893_ff <= lut_1893_out;
            end
        end
        
        assign out_data[1893] = lut_1893_ff;
    end
    else begin : no_ff_1893
        assign out_data[1893] = lut_1893_out;
    end
    endgenerate
    
    
    
    // LUT : 1894
    wire [63:0] lut_1894_table = 64'b1111000000000010111111111111110011111100110011001111111111000100;
    wire [5:0] lut_1894_select = {
                             in_data[400],
                             in_data[658],
                             in_data[488],
                             in_data[377],
                             in_data[583],
                             in_data[765]};
    
    wire lut_1894_out = lut_1894_table[lut_1894_select];
    
    generate
    if ( USE_REG ) begin : ff_1894
        reg   lut_1894_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1894_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1894_ff <= lut_1894_out;
            end
        end
        
        assign out_data[1894] = lut_1894_ff;
    end
    else begin : no_ff_1894
        assign out_data[1894] = lut_1894_out;
    end
    endgenerate
    
    
    
    // LUT : 1895
    wire [63:0] lut_1895_table = 64'b0000000000000000111111111111111100000000000000001110101011111010;
    wire [5:0] lut_1895_select = {
                             in_data[199],
                             in_data[651],
                             in_data[217],
                             in_data[290],
                             in_data[2],
                             in_data[64]};
    
    wire lut_1895_out = lut_1895_table[lut_1895_select];
    
    generate
    if ( USE_REG ) begin : ff_1895
        reg   lut_1895_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1895_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1895_ff <= lut_1895_out;
            end
        end
        
        assign out_data[1895] = lut_1895_ff;
    end
    else begin : no_ff_1895
        assign out_data[1895] = lut_1895_out;
    end
    endgenerate
    
    
    
    // LUT : 1896
    wire [63:0] lut_1896_table = 64'b0000000011001111000000001100110100000000110011110000000011001101;
    wire [5:0] lut_1896_select = {
                             in_data[778],
                             in_data[137],
                             in_data[319],
                             in_data[677],
                             in_data[288],
                             in_data[86]};
    
    wire lut_1896_out = lut_1896_table[lut_1896_select];
    
    generate
    if ( USE_REG ) begin : ff_1896
        reg   lut_1896_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1896_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1896_ff <= lut_1896_out;
            end
        end
        
        assign out_data[1896] = lut_1896_ff;
    end
    else begin : no_ff_1896
        assign out_data[1896] = lut_1896_out;
    end
    endgenerate
    
    
    
    // LUT : 1897
    wire [63:0] lut_1897_table = 64'b1011111100101011001010110010001110111111001010110011101100100011;
    wire [5:0] lut_1897_select = {
                             in_data[780],
                             in_data[160],
                             in_data[648],
                             in_data[345],
                             in_data[694],
                             in_data[147]};
    
    wire lut_1897_out = lut_1897_table[lut_1897_select];
    
    generate
    if ( USE_REG ) begin : ff_1897
        reg   lut_1897_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1897_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1897_ff <= lut_1897_out;
            end
        end
        
        assign out_data[1897] = lut_1897_ff;
    end
    else begin : no_ff_1897
        assign out_data[1897] = lut_1897_out;
    end
    endgenerate
    
    
    
    // LUT : 1898
    wire [63:0] lut_1898_table = 64'b0011001100110011001100110011001100100010001000100010001000100010;
    wire [5:0] lut_1898_select = {
                             in_data[387],
                             in_data[60],
                             in_data[112],
                             in_data[753],
                             in_data[266],
                             in_data[494]};
    
    wire lut_1898_out = lut_1898_table[lut_1898_select];
    
    generate
    if ( USE_REG ) begin : ff_1898
        reg   lut_1898_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1898_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1898_ff <= lut_1898_out;
            end
        end
        
        assign out_data[1898] = lut_1898_ff;
    end
    else begin : no_ff_1898
        assign out_data[1898] = lut_1898_out;
    end
    endgenerate
    
    
    
    // LUT : 1899
    wire [63:0] lut_1899_table = 64'b1111111111111111000000010000000011111111111111110000000100000000;
    wire [5:0] lut_1899_select = {
                             in_data[62],
                             in_data[153],
                             in_data[268],
                             in_data[361],
                             in_data[716],
                             in_data[163]};
    
    wire lut_1899_out = lut_1899_table[lut_1899_select];
    
    generate
    if ( USE_REG ) begin : ff_1899
        reg   lut_1899_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1899_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1899_ff <= lut_1899_out;
            end
        end
        
        assign out_data[1899] = lut_1899_ff;
    end
    else begin : no_ff_1899
        assign out_data[1899] = lut_1899_out;
    end
    endgenerate
    
    
    
    // LUT : 1900
    wire [63:0] lut_1900_table = 64'b0000010100000001001101110011011100000001000000010001011100010111;
    wire [5:0] lut_1900_select = {
                             in_data[622],
                             in_data[292],
                             in_data[613],
                             in_data[276],
                             in_data[510],
                             in_data[242]};
    
    wire lut_1900_out = lut_1900_table[lut_1900_select];
    
    generate
    if ( USE_REG ) begin : ff_1900
        reg   lut_1900_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1900_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1900_ff <= lut_1900_out;
            end
        end
        
        assign out_data[1900] = lut_1900_ff;
    end
    else begin : no_ff_1900
        assign out_data[1900] = lut_1900_out;
    end
    endgenerate
    
    
    
    // LUT : 1901
    wire [63:0] lut_1901_table = 64'b0000010100001111110011010000111111001100110011001100110011001100;
    wire [5:0] lut_1901_select = {
                             in_data[182],
                             in_data[5],
                             in_data[484],
                             in_data[425],
                             in_data[126],
                             in_data[702]};
    
    wire lut_1901_out = lut_1901_table[lut_1901_select];
    
    generate
    if ( USE_REG ) begin : ff_1901
        reg   lut_1901_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1901_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1901_ff <= lut_1901_out;
            end
        end
        
        assign out_data[1901] = lut_1901_ff;
    end
    else begin : no_ff_1901
        assign out_data[1901] = lut_1901_out;
    end
    endgenerate
    
    
    
    // LUT : 1902
    wire [63:0] lut_1902_table = 64'b0000000000001111000000110000101100000000000000000000000100000011;
    wire [5:0] lut_1902_select = {
                             in_data[526],
                             in_data[598],
                             in_data[216],
                             in_data[258],
                             in_data[710],
                             in_data[637]};
    
    wire lut_1902_out = lut_1902_table[lut_1902_select];
    
    generate
    if ( USE_REG ) begin : ff_1902
        reg   lut_1902_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1902_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1902_ff <= lut_1902_out;
            end
        end
        
        assign out_data[1902] = lut_1902_ff;
    end
    else begin : no_ff_1902
        assign out_data[1902] = lut_1902_out;
    end
    endgenerate
    
    
    
    // LUT : 1903
    wire [63:0] lut_1903_table = 64'b1100110011001100110011001100110011111110111111101111111011111110;
    wire [5:0] lut_1903_select = {
                             in_data[373],
                             in_data[569],
                             in_data[531],
                             in_data[282],
                             in_data[384],
                             in_data[751]};
    
    wire lut_1903_out = lut_1903_table[lut_1903_select];
    
    generate
    if ( USE_REG ) begin : ff_1903
        reg   lut_1903_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1903_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1903_ff <= lut_1903_out;
            end
        end
        
        assign out_data[1903] = lut_1903_ff;
    end
    else begin : no_ff_1903
        assign out_data[1903] = lut_1903_out;
    end
    endgenerate
    
    
    
    // LUT : 1904
    wire [63:0] lut_1904_table = 64'b1111111111111111111111111111111111111111111111110000000000000000;
    wire [5:0] lut_1904_select = {
                             in_data[423],
                             in_data[293],
                             in_data[9],
                             in_data[117],
                             in_data[135],
                             in_data[777]};
    
    wire lut_1904_out = lut_1904_table[lut_1904_select];
    
    generate
    if ( USE_REG ) begin : ff_1904
        reg   lut_1904_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1904_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1904_ff <= lut_1904_out;
            end
        end
        
        assign out_data[1904] = lut_1904_ff;
    end
    else begin : no_ff_1904
        assign out_data[1904] = lut_1904_out;
    end
    endgenerate
    
    
    
    // LUT : 1905
    wire [63:0] lut_1905_table = 64'b1111111100110011111111110011000011111111001100111111111100110000;
    wire [5:0] lut_1905_select = {
                             in_data[586],
                             in_data[545],
                             in_data[321],
                             in_data[536],
                             in_data[357],
                             in_data[417]};
    
    wire lut_1905_out = lut_1905_table[lut_1905_select];
    
    generate
    if ( USE_REG ) begin : ff_1905
        reg   lut_1905_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1905_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1905_ff <= lut_1905_out;
            end
        end
        
        assign out_data[1905] = lut_1905_ff;
    end
    else begin : no_ff_1905
        assign out_data[1905] = lut_1905_out;
    end
    endgenerate
    
    
    
    // LUT : 1906
    wire [63:0] lut_1906_table = 64'b0000000000000000000000000000000000000000000000000000000001111111;
    wire [5:0] lut_1906_select = {
                             in_data[584],
                             in_data[155],
                             in_data[553],
                             in_data[29],
                             in_data[414],
                             in_data[775]};
    
    wire lut_1906_out = lut_1906_table[lut_1906_select];
    
    generate
    if ( USE_REG ) begin : ff_1906
        reg   lut_1906_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1906_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1906_ff <= lut_1906_out;
            end
        end
        
        assign out_data[1906] = lut_1906_ff;
    end
    else begin : no_ff_1906
        assign out_data[1906] = lut_1906_out;
    end
    endgenerate
    
    
    
    // LUT : 1907
    wire [63:0] lut_1907_table = 64'b0000000000000000000000000000000011101111111111111110111011111111;
    wire [5:0] lut_1907_select = {
                             in_data[407],
                             in_data[410],
                             in_data[680],
                             in_data[615],
                             in_data[76],
                             in_data[238]};
    
    wire lut_1907_out = lut_1907_table[lut_1907_select];
    
    generate
    if ( USE_REG ) begin : ff_1907
        reg   lut_1907_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1907_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1907_ff <= lut_1907_out;
            end
        end
        
        assign out_data[1907] = lut_1907_ff;
    end
    else begin : no_ff_1907
        assign out_data[1907] = lut_1907_out;
    end
    endgenerate
    
    
    
    // LUT : 1908
    wire [63:0] lut_1908_table = 64'b0011001100110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1908_select = {
                             in_data[750],
                             in_data[587],
                             in_data[684],
                             in_data[104],
                             in_data[329],
                             in_data[486]};
    
    wire lut_1908_out = lut_1908_table[lut_1908_select];
    
    generate
    if ( USE_REG ) begin : ff_1908
        reg   lut_1908_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1908_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1908_ff <= lut_1908_out;
            end
        end
        
        assign out_data[1908] = lut_1908_ff;
    end
    else begin : no_ff_1908
        assign out_data[1908] = lut_1908_out;
    end
    endgenerate
    
    
    
    // LUT : 1909
    wire [63:0] lut_1909_table = 64'b0000000000000000010101010000000011111111111111111111111111111010;
    wire [5:0] lut_1909_select = {
                             in_data[404],
                             in_data[316],
                             in_data[228],
                             in_data[512],
                             in_data[390],
                             in_data[455]};
    
    wire lut_1909_out = lut_1909_table[lut_1909_select];
    
    generate
    if ( USE_REG ) begin : ff_1909
        reg   lut_1909_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1909_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1909_ff <= lut_1909_out;
            end
        end
        
        assign out_data[1909] = lut_1909_ff;
    end
    else begin : no_ff_1909
        assign out_data[1909] = lut_1909_out;
    end
    endgenerate
    
    
    
    // LUT : 1910
    wire [63:0] lut_1910_table = 64'b1111111111111111001000100010001011111111111111111010001010101010;
    wire [5:0] lut_1910_select = {
                             in_data[362],
                             in_data[131],
                             in_data[767],
                             in_data[39],
                             in_data[463],
                             in_data[237]};
    
    wire lut_1910_out = lut_1910_table[lut_1910_select];
    
    generate
    if ( USE_REG ) begin : ff_1910
        reg   lut_1910_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1910_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1910_ff <= lut_1910_out;
            end
        end
        
        assign out_data[1910] = lut_1910_ff;
    end
    else begin : no_ff_1910
        assign out_data[1910] = lut_1910_out;
    end
    endgenerate
    
    
    
    // LUT : 1911
    wire [63:0] lut_1911_table = 64'b0000000000000000111111100100010000000000000000001111111101010101;
    wire [5:0] lut_1911_select = {
                             in_data[310],
                             in_data[256],
                             in_data[466],
                             in_data[421],
                             in_data[307],
                             in_data[630]};
    
    wire lut_1911_out = lut_1911_table[lut_1911_select];
    
    generate
    if ( USE_REG ) begin : ff_1911
        reg   lut_1911_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1911_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1911_ff <= lut_1911_out;
            end
        end
        
        assign out_data[1911] = lut_1911_ff;
    end
    else begin : no_ff_1911
        assign out_data[1911] = lut_1911_out;
    end
    endgenerate
    
    
    
    // LUT : 1912
    wire [63:0] lut_1912_table = 64'b0000000000000000000000000000000011010101110111011101110111011101;
    wire [5:0] lut_1912_select = {
                             in_data[356],
                             in_data[749],
                             in_data[641],
                             in_data[193],
                             in_data[578],
                             in_data[551]};
    
    wire lut_1912_out = lut_1912_table[lut_1912_select];
    
    generate
    if ( USE_REG ) begin : ff_1912
        reg   lut_1912_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1912_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1912_ff <= lut_1912_out;
            end
        end
        
        assign out_data[1912] = lut_1912_ff;
    end
    else begin : no_ff_1912
        assign out_data[1912] = lut_1912_out;
    end
    endgenerate
    
    
    
    // LUT : 1913
    wire [63:0] lut_1913_table = 64'b0000000000000000000000000000000000111011001110110011001000111010;
    wire [5:0] lut_1913_select = {
                             in_data[564],
                             in_data[226],
                             in_data[79],
                             in_data[313],
                             in_data[603],
                             in_data[408]};
    
    wire lut_1913_out = lut_1913_table[lut_1913_select];
    
    generate
    if ( USE_REG ) begin : ff_1913
        reg   lut_1913_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1913_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1913_ff <= lut_1913_out;
            end
        end
        
        assign out_data[1913] = lut_1913_ff;
    end
    else begin : no_ff_1913
        assign out_data[1913] = lut_1913_out;
    end
    endgenerate
    
    
    
    // LUT : 1914
    wire [63:0] lut_1914_table = 64'b0000000000000000000000000000000010100000100000001110111111101111;
    wire [5:0] lut_1914_select = {
                             in_data[580],
                             in_data[180],
                             in_data[755],
                             in_data[257],
                             in_data[109],
                             in_data[415]};
    
    wire lut_1914_out = lut_1914_table[lut_1914_select];
    
    generate
    if ( USE_REG ) begin : ff_1914
        reg   lut_1914_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1914_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1914_ff <= lut_1914_out;
            end
        end
        
        assign out_data[1914] = lut_1914_ff;
    end
    else begin : no_ff_1914
        assign out_data[1914] = lut_1914_out;
    end
    endgenerate
    
    
    
    // LUT : 1915
    wire [63:0] lut_1915_table = 64'b1101110011011100110111001101110011011100110111001101110011011100;
    wire [5:0] lut_1915_select = {
                             in_data[448],
                             in_data[8],
                             in_data[166],
                             in_data[100],
                             in_data[544],
                             in_data[96]};
    
    wire lut_1915_out = lut_1915_table[lut_1915_select];
    
    generate
    if ( USE_REG ) begin : ff_1915
        reg   lut_1915_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1915_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1915_ff <= lut_1915_out;
            end
        end
        
        assign out_data[1915] = lut_1915_ff;
    end
    else begin : no_ff_1915
        assign out_data[1915] = lut_1915_out;
    end
    endgenerate
    
    
    
    // LUT : 1916
    wire [63:0] lut_1916_table = 64'b0000000000000000000000000000000100000000000101010000000000000101;
    wire [5:0] lut_1916_select = {
                             in_data[469],
                             in_data[733],
                             in_data[118],
                             in_data[382],
                             in_data[84],
                             in_data[682]};
    
    wire lut_1916_out = lut_1916_table[lut_1916_select];
    
    generate
    if ( USE_REG ) begin : ff_1916
        reg   lut_1916_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1916_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1916_ff <= lut_1916_out;
            end
        end
        
        assign out_data[1916] = lut_1916_ff;
    end
    else begin : no_ff_1916
        assign out_data[1916] = lut_1916_out;
    end
    endgenerate
    
    
    
    // LUT : 1917
    wire [63:0] lut_1917_table = 64'b1111111111111111111111111111111111101110111011101100110011001110;
    wire [5:0] lut_1917_select = {
                             in_data[205],
                             in_data[41],
                             in_data[12],
                             in_data[614],
                             in_data[600],
                             in_data[507]};
    
    wire lut_1917_out = lut_1917_table[lut_1917_select];
    
    generate
    if ( USE_REG ) begin : ff_1917
        reg   lut_1917_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1917_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1917_ff <= lut_1917_out;
            end
        end
        
        assign out_data[1917] = lut_1917_ff;
    end
    else begin : no_ff_1917
        assign out_data[1917] = lut_1917_out;
    end
    endgenerate
    
    
    
    // LUT : 1918
    wire [63:0] lut_1918_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_1918_select = {
                             in_data[559],
                             in_data[263],
                             in_data[418],
                             in_data[103],
                             in_data[17],
                             in_data[291]};
    
    wire lut_1918_out = lut_1918_table[lut_1918_select];
    
    generate
    if ( USE_REG ) begin : ff_1918
        reg   lut_1918_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1918_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1918_ff <= lut_1918_out;
            end
        end
        
        assign out_data[1918] = lut_1918_ff;
    end
    else begin : no_ff_1918
        assign out_data[1918] = lut_1918_out;
    end
    endgenerate
    
    
    
    // LUT : 1919
    wire [63:0] lut_1919_table = 64'b0100010000000000000000000000000011101110010101011010111011111111;
    wire [5:0] lut_1919_select = {
                             in_data[323],
                             in_data[245],
                             in_data[579],
                             in_data[768],
                             in_data[368],
                             in_data[546]};
    
    wire lut_1919_out = lut_1919_table[lut_1919_select];
    
    generate
    if ( USE_REG ) begin : ff_1919
        reg   lut_1919_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1919_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1919_ff <= lut_1919_out;
            end
        end
        
        assign out_data[1919] = lut_1919_ff;
    end
    else begin : no_ff_1919
        assign out_data[1919] = lut_1919_out;
    end
    endgenerate
    
    
    
    // LUT : 1920
    wire [63:0] lut_1920_table = 64'b0101000100010000010101010101000101010001010100000101010101010001;
    wire [5:0] lut_1920_select = {
                             in_data[670],
                             in_data[249],
                             in_data[209],
                             in_data[443],
                             in_data[746],
                             in_data[628]};
    
    wire lut_1920_out = lut_1920_table[lut_1920_select];
    
    generate
    if ( USE_REG ) begin : ff_1920
        reg   lut_1920_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1920_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1920_ff <= lut_1920_out;
            end
        end
        
        assign out_data[1920] = lut_1920_ff;
    end
    else begin : no_ff_1920
        assign out_data[1920] = lut_1920_out;
    end
    endgenerate
    
    
    
    // LUT : 1921
    wire [63:0] lut_1921_table = 64'b1111000011110000111100001111000011110000111100001111000011110101;
    wire [5:0] lut_1921_select = {
                             in_data[239],
                             in_data[688],
                             in_data[349],
                             in_data[270],
                             in_data[697],
                             in_data[68]};
    
    wire lut_1921_out = lut_1921_table[lut_1921_select];
    
    generate
    if ( USE_REG ) begin : ff_1921
        reg   lut_1921_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1921_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1921_ff <= lut_1921_out;
            end
        end
        
        assign out_data[1921] = lut_1921_ff;
    end
    else begin : no_ff_1921
        assign out_data[1921] = lut_1921_out;
    end
    endgenerate
    
    
    
    // LUT : 1922
    wire [63:0] lut_1922_table = 64'b0000010100000101000001010000010100000101000001010000010100000101;
    wire [5:0] lut_1922_select = {
                             in_data[4],
                             in_data[644],
                             in_data[491],
                             in_data[480],
                             in_data[392],
                             in_data[490]};
    
    wire lut_1922_out = lut_1922_table[lut_1922_select];
    
    generate
    if ( USE_REG ) begin : ff_1922
        reg   lut_1922_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1922_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1922_ff <= lut_1922_out;
            end
        end
        
        assign out_data[1922] = lut_1922_ff;
    end
    else begin : no_ff_1922
        assign out_data[1922] = lut_1922_out;
    end
    endgenerate
    
    
    
    // LUT : 1923
    wire [63:0] lut_1923_table = 64'b0000000011110111000000000101000100010001000100010001000100010001;
    wire [5:0] lut_1923_select = {
                             in_data[208],
                             in_data[73],
                             in_data[689],
                             in_data[704],
                             in_data[568],
                             in_data[713]};
    
    wire lut_1923_out = lut_1923_table[lut_1923_select];
    
    generate
    if ( USE_REG ) begin : ff_1923
        reg   lut_1923_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1923_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1923_ff <= lut_1923_out;
            end
        end
        
        assign out_data[1923] = lut_1923_ff;
    end
    else begin : no_ff_1923
        assign out_data[1923] = lut_1923_out;
    end
    endgenerate
    
    
    
    // LUT : 1924
    wire [63:0] lut_1924_table = 64'b0000000000000000000000000000000000000000010111110000000000001111;
    wire [5:0] lut_1924_select = {
                             in_data[550],
                             in_data[35],
                             in_data[250],
                             in_data[576],
                             in_data[57],
                             in_data[114]};
    
    wire lut_1924_out = lut_1924_table[lut_1924_select];
    
    generate
    if ( USE_REG ) begin : ff_1924
        reg   lut_1924_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1924_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1924_ff <= lut_1924_out;
            end
        end
        
        assign out_data[1924] = lut_1924_ff;
    end
    else begin : no_ff_1924
        assign out_data[1924] = lut_1924_out;
    end
    endgenerate
    
    
    
    // LUT : 1925
    wire [63:0] lut_1925_table = 64'b1111111111111111111111111111111100000000001100110011000000110010;
    wire [5:0] lut_1925_select = {
                             in_data[571],
                             in_data[364],
                             in_data[566],
                             in_data[20],
                             in_data[438],
                             in_data[34]};
    
    wire lut_1925_out = lut_1925_table[lut_1925_select];
    
    generate
    if ( USE_REG ) begin : ff_1925
        reg   lut_1925_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1925_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1925_ff <= lut_1925_out;
            end
        end
        
        assign out_data[1925] = lut_1925_ff;
    end
    else begin : no_ff_1925
        assign out_data[1925] = lut_1925_out;
    end
    endgenerate
    
    
    
    // LUT : 1926
    wire [63:0] lut_1926_table = 64'b0000000100000011000000110000001100110011001100110011101100110011;
    wire [5:0] lut_1926_select = {
                             in_data[611],
                             in_data[640],
                             in_data[3],
                             in_data[264],
                             in_data[431],
                             in_data[14]};
    
    wire lut_1926_out = lut_1926_table[lut_1926_select];
    
    generate
    if ( USE_REG ) begin : ff_1926
        reg   lut_1926_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1926_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1926_ff <= lut_1926_out;
            end
        end
        
        assign out_data[1926] = lut_1926_ff;
    end
    else begin : no_ff_1926
        assign out_data[1926] = lut_1926_out;
    end
    endgenerate
    
    
    
    // LUT : 1927
    wire [63:0] lut_1927_table = 64'b0000000010001010000000001000100011111111111111111111111011111111;
    wire [5:0] lut_1927_select = {
                             in_data[157],
                             in_data[783],
                             in_data[317],
                             in_data[344],
                             in_data[66],
                             in_data[721]};
    
    wire lut_1927_out = lut_1927_table[lut_1927_select];
    
    generate
    if ( USE_REG ) begin : ff_1927
        reg   lut_1927_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1927_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1927_ff <= lut_1927_out;
            end
        end
        
        assign out_data[1927] = lut_1927_ff;
    end
    else begin : no_ff_1927
        assign out_data[1927] = lut_1927_out;
    end
    endgenerate
    
    
    
    // LUT : 1928
    wire [63:0] lut_1928_table = 64'b0100111101001111000001000000010011001111110011110000110100001100;
    wire [5:0] lut_1928_select = {
                             in_data[394],
                             in_data[40],
                             in_data[726],
                             in_data[719],
                             in_data[119],
                             in_data[143]};
    
    wire lut_1928_out = lut_1928_table[lut_1928_select];
    
    generate
    if ( USE_REG ) begin : ff_1928
        reg   lut_1928_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1928_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1928_ff <= lut_1928_out;
            end
        end
        
        assign out_data[1928] = lut_1928_ff;
    end
    else begin : no_ff_1928
        assign out_data[1928] = lut_1928_out;
    end
    endgenerate
    
    
    
    // LUT : 1929
    wire [63:0] lut_1929_table = 64'b1111111111111111000000001111111111111111111111110000000011111111;
    wire [5:0] lut_1929_select = {
                             in_data[758],
                             in_data[683],
                             in_data[325],
                             in_data[592],
                             in_data[223],
                             in_data[27]};
    
    wire lut_1929_out = lut_1929_table[lut_1929_select];
    
    generate
    if ( USE_REG ) begin : ff_1929
        reg   lut_1929_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1929_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1929_ff <= lut_1929_out;
            end
        end
        
        assign out_data[1929] = lut_1929_ff;
    end
    else begin : no_ff_1929
        assign out_data[1929] = lut_1929_out;
    end
    endgenerate
    
    
    
    // LUT : 1930
    wire [63:0] lut_1930_table = 64'b1111111111111111010000000101010111111111111111110101000101010101;
    wire [5:0] lut_1930_select = {
                             in_data[90],
                             in_data[623],
                             in_data[675],
                             in_data[31],
                             in_data[724],
                             in_data[235]};
    
    wire lut_1930_out = lut_1930_table[lut_1930_select];
    
    generate
    if ( USE_REG ) begin : ff_1930
        reg   lut_1930_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1930_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1930_ff <= lut_1930_out;
            end
        end
        
        assign out_data[1930] = lut_1930_ff;
    end
    else begin : no_ff_1930
        assign out_data[1930] = lut_1930_out;
    end
    endgenerate
    
    
    
    // LUT : 1931
    wire [63:0] lut_1931_table = 64'b1111111111111111111101011111010100001010000010100000000000000000;
    wire [5:0] lut_1931_select = {
                             in_data[570],
                             in_data[244],
                             in_data[37],
                             in_data[492],
                             in_data[504],
                             in_data[246]};
    
    wire lut_1931_out = lut_1931_table[lut_1931_select];
    
    generate
    if ( USE_REG ) begin : ff_1931
        reg   lut_1931_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1931_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1931_ff <= lut_1931_out;
            end
        end
        
        assign out_data[1931] = lut_1931_ff;
    end
    else begin : no_ff_1931
        assign out_data[1931] = lut_1931_out;
    end
    endgenerate
    
    
    
    // LUT : 1932
    wire [63:0] lut_1932_table = 64'b1111010111110101111101011111010111110101111101011111010111110101;
    wire [5:0] lut_1932_select = {
                             in_data[252],
                             in_data[141],
                             in_data[138],
                             in_data[609],
                             in_data[478],
                             in_data[409]};
    
    wire lut_1932_out = lut_1932_table[lut_1932_select];
    
    generate
    if ( USE_REG ) begin : ff_1932
        reg   lut_1932_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1932_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1932_ff <= lut_1932_out;
            end
        end
        
        assign out_data[1932] = lut_1932_ff;
    end
    else begin : no_ff_1932
        assign out_data[1932] = lut_1932_out;
    end
    endgenerate
    
    
    
    // LUT : 1933
    wire [63:0] lut_1933_table = 64'b1000100010001000110010011100110110001000100010001100100111011001;
    wire [5:0] lut_1933_select = {
                             in_data[47],
                             in_data[433],
                             in_data[65],
                             in_data[520],
                             in_data[625],
                             in_data[572]};
    
    wire lut_1933_out = lut_1933_table[lut_1933_select];
    
    generate
    if ( USE_REG ) begin : ff_1933
        reg   lut_1933_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1933_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1933_ff <= lut_1933_out;
            end
        end
        
        assign out_data[1933] = lut_1933_ff;
    end
    else begin : no_ff_1933
        assign out_data[1933] = lut_1933_out;
    end
    endgenerate
    
    
    
    // LUT : 1934
    wire [63:0] lut_1934_table = 64'b0000000000000000010101010101010100000000000000000101010101010101;
    wire [5:0] lut_1934_select = {
                             in_data[560],
                             in_data[332],
                             in_data[111],
                             in_data[142],
                             in_data[712],
                             in_data[183]};
    
    wire lut_1934_out = lut_1934_table[lut_1934_select];
    
    generate
    if ( USE_REG ) begin : ff_1934
        reg   lut_1934_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1934_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1934_ff <= lut_1934_out;
            end
        end
        
        assign out_data[1934] = lut_1934_ff;
    end
    else begin : no_ff_1934
        assign out_data[1934] = lut_1934_out;
    end
    endgenerate
    
    
    
    // LUT : 1935
    wire [63:0] lut_1935_table = 64'b1111111111111111111111111010101011111111111111111111111110101010;
    wire [5:0] lut_1935_select = {
                             in_data[43],
                             in_data[539],
                             in_data[101],
                             in_data[365],
                             in_data[279],
                             in_data[98]};
    
    wire lut_1935_out = lut_1935_table[lut_1935_select];
    
    generate
    if ( USE_REG ) begin : ff_1935
        reg   lut_1935_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1935_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1935_ff <= lut_1935_out;
            end
        end
        
        assign out_data[1935] = lut_1935_ff;
    end
    else begin : no_ff_1935
        assign out_data[1935] = lut_1935_out;
    end
    endgenerate
    
    
    
    // LUT : 1936
    wire [63:0] lut_1936_table = 64'b0000111100001010000111110000111100001111000010100001111100001111;
    wire [5:0] lut_1936_select = {
                             in_data[24],
                             in_data[735],
                             in_data[585],
                             in_data[573],
                             in_data[371],
                             in_data[496]};
    
    wire lut_1936_out = lut_1936_table[lut_1936_select];
    
    generate
    if ( USE_REG ) begin : ff_1936
        reg   lut_1936_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1936_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1936_ff <= lut_1936_out;
            end
        end
        
        assign out_data[1936] = lut_1936_ff;
    end
    else begin : no_ff_1936
        assign out_data[1936] = lut_1936_out;
    end
    endgenerate
    
    
    
    // LUT : 1937
    wire [63:0] lut_1937_table = 64'b0000000011111111000000000000000000000000111111110000000000000000;
    wire [5:0] lut_1937_select = {
                             in_data[30],
                             in_data[212],
                             in_data[518],
                             in_data[234],
                             in_data[80],
                             in_data[343]};
    
    wire lut_1937_out = lut_1937_table[lut_1937_select];
    
    generate
    if ( USE_REG ) begin : ff_1937
        reg   lut_1937_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1937_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1937_ff <= lut_1937_out;
            end
        end
        
        assign out_data[1937] = lut_1937_ff;
    end
    else begin : no_ff_1937
        assign out_data[1937] = lut_1937_out;
    end
    endgenerate
    
    
    
    // LUT : 1938
    wire [63:0] lut_1938_table = 64'b1111111100000011111111111100001111001110000000001111111100000000;
    wire [5:0] lut_1938_select = {
                             in_data[174],
                             in_data[772],
                             in_data[483],
                             in_data[633],
                             in_data[457],
                             in_data[393]};
    
    wire lut_1938_out = lut_1938_table[lut_1938_select];
    
    generate
    if ( USE_REG ) begin : ff_1938
        reg   lut_1938_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1938_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1938_ff <= lut_1938_out;
            end
        end
        
        assign out_data[1938] = lut_1938_ff;
    end
    else begin : no_ff_1938
        assign out_data[1938] = lut_1938_out;
    end
    endgenerate
    
    
    
    // LUT : 1939
    wire [63:0] lut_1939_table = 64'b1110111111111111000011110000111100001111010011110000000000000000;
    wire [5:0] lut_1939_select = {
                             in_data[656],
                             in_data[331],
                             in_data[695],
                             in_data[717],
                             in_data[419],
                             in_data[336]};
    
    wire lut_1939_out = lut_1939_table[lut_1939_select];
    
    generate
    if ( USE_REG ) begin : ff_1939
        reg   lut_1939_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1939_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1939_ff <= lut_1939_out;
            end
        end
        
        assign out_data[1939] = lut_1939_ff;
    end
    else begin : no_ff_1939
        assign out_data[1939] = lut_1939_out;
    end
    endgenerate
    
    
    
    // LUT : 1940
    wire [63:0] lut_1940_table = 64'b1111111111111111111111111111111111111111101011110000101100000000;
    wire [5:0] lut_1940_select = {
                             in_data[127],
                             in_data[399],
                             in_data[720],
                             in_data[403],
                             in_data[781],
                             in_data[445]};
    
    wire lut_1940_out = lut_1940_table[lut_1940_select];
    
    generate
    if ( USE_REG ) begin : ff_1940
        reg   lut_1940_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1940_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1940_ff <= lut_1940_out;
            end
        end
        
        assign out_data[1940] = lut_1940_ff;
    end
    else begin : no_ff_1940
        assign out_data[1940] = lut_1940_out;
    end
    endgenerate
    
    
    
    // LUT : 1941
    wire [63:0] lut_1941_table = 64'b0010111100100010000000100000000011111111111111110010001100100011;
    wire [5:0] lut_1941_select = {
                             in_data[556],
                             in_data[397],
                             in_data[391],
                             in_data[164],
                             in_data[185],
                             in_data[691]};
    
    wire lut_1941_out = lut_1941_table[lut_1941_select];
    
    generate
    if ( USE_REG ) begin : ff_1941
        reg   lut_1941_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1941_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1941_ff <= lut_1941_out;
            end
        end
        
        assign out_data[1941] = lut_1941_ff;
    end
    else begin : no_ff_1941
        assign out_data[1941] = lut_1941_out;
    end
    endgenerate
    
    
    
    // LUT : 1942
    wire [63:0] lut_1942_table = 64'b0000000000000000000010100000101000000000000000000000101010101010;
    wire [5:0] lut_1942_select = {
                             in_data[275],
                             in_data[621],
                             in_data[561],
                             in_data[348],
                             in_data[59],
                             in_data[437]};
    
    wire lut_1942_out = lut_1942_table[lut_1942_select];
    
    generate
    if ( USE_REG ) begin : ff_1942
        reg   lut_1942_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1942_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1942_ff <= lut_1942_out;
            end
        end
        
        assign out_data[1942] = lut_1942_ff;
    end
    else begin : no_ff_1942
        assign out_data[1942] = lut_1942_out;
    end
    endgenerate
    
    
    
    // LUT : 1943
    wire [63:0] lut_1943_table = 64'b0011000011111100000000001100110011110010111111110000000011111100;
    wire [5:0] lut_1943_select = {
                             in_data[312],
                             in_data[685],
                             in_data[102],
                             in_data[555],
                             in_data[629],
                             in_data[18]};
    
    wire lut_1943_out = lut_1943_table[lut_1943_select];
    
    generate
    if ( USE_REG ) begin : ff_1943
        reg   lut_1943_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1943_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1943_ff <= lut_1943_out;
            end
        end
        
        assign out_data[1943] = lut_1943_ff;
    end
    else begin : no_ff_1943
        assign out_data[1943] = lut_1943_out;
    end
    endgenerate
    
    
    
    // LUT : 1944
    wire [63:0] lut_1944_table = 64'b1111101111111011001100110011001100000000000000001111111100110011;
    wire [5:0] lut_1944_select = {
                             in_data[542],
                             in_data[459],
                             in_data[302],
                             in_data[0],
                             in_data[233],
                             in_data[477]};
    
    wire lut_1944_out = lut_1944_table[lut_1944_select];
    
    generate
    if ( USE_REG ) begin : ff_1944
        reg   lut_1944_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1944_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1944_ff <= lut_1944_out;
            end
        end
        
        assign out_data[1944] = lut_1944_ff;
    end
    else begin : no_ff_1944
        assign out_data[1944] = lut_1944_out;
    end
    endgenerate
    
    
    
    // LUT : 1945
    wire [63:0] lut_1945_table = 64'b0000010001000101000001000100010111001101110111011100110111011101;
    wire [5:0] lut_1945_select = {
                             in_data[411],
                             in_data[643],
                             in_data[740],
                             in_data[426],
                             in_data[678],
                             in_data[517]};
    
    wire lut_1945_out = lut_1945_table[lut_1945_select];
    
    generate
    if ( USE_REG ) begin : ff_1945
        reg   lut_1945_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1945_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1945_ff <= lut_1945_out;
            end
        end
        
        assign out_data[1945] = lut_1945_ff;
    end
    else begin : no_ff_1945
        assign out_data[1945] = lut_1945_out;
    end
    endgenerate
    
    
    
    // LUT : 1946
    wire [63:0] lut_1946_table = 64'b1111000011110000111100001111000011111100111110001111110011111100;
    wire [5:0] lut_1946_select = {
                             in_data[240],
                             in_data[725],
                             in_data[13],
                             in_data[210],
                             in_data[436],
                             in_data[225]};
    
    wire lut_1946_out = lut_1946_table[lut_1946_select];
    
    generate
    if ( USE_REG ) begin : ff_1946
        reg   lut_1946_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1946_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1946_ff <= lut_1946_out;
            end
        end
        
        assign out_data[1946] = lut_1946_ff;
    end
    else begin : no_ff_1946
        assign out_data[1946] = lut_1946_out;
    end
    endgenerate
    
    
    
    // LUT : 1947
    wire [63:0] lut_1947_table = 64'b0010000011001100001000001100110100110100110011010011010011001101;
    wire [5:0] lut_1947_select = {
                             in_data[110],
                             in_data[698],
                             in_data[430],
                             in_data[158],
                             in_data[267],
                             in_data[515]};
    
    wire lut_1947_out = lut_1947_table[lut_1947_select];
    
    generate
    if ( USE_REG ) begin : ff_1947
        reg   lut_1947_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1947_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1947_ff <= lut_1947_out;
            end
        end
        
        assign out_data[1947] = lut_1947_ff;
    end
    else begin : no_ff_1947
        assign out_data[1947] = lut_1947_out;
    end
    endgenerate
    
    
    
    // LUT : 1948
    wire [63:0] lut_1948_table = 64'b1111100011111111000000001100110011111000111111110000000011001100;
    wire [5:0] lut_1948_select = {
                             in_data[779],
                             in_data[528],
                             in_data[333],
                             in_data[524],
                             in_data[485],
                             in_data[475]};
    
    wire lut_1948_out = lut_1948_table[lut_1948_select];
    
    generate
    if ( USE_REG ) begin : ff_1948
        reg   lut_1948_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1948_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1948_ff <= lut_1948_out;
            end
        end
        
        assign out_data[1948] = lut_1948_ff;
    end
    else begin : no_ff_1948
        assign out_data[1948] = lut_1948_out;
    end
    endgenerate
    
    
    
    // LUT : 1949
    wire [63:0] lut_1949_table = 64'b1100111111001110110011111100111000000010000011100000011000001110;
    wire [5:0] lut_1949_select = {
                             in_data[346],
                             in_data[83],
                             in_data[442],
                             in_data[359],
                             in_data[606],
                             in_data[204]};
    
    wire lut_1949_out = lut_1949_table[lut_1949_select];
    
    generate
    if ( USE_REG ) begin : ff_1949
        reg   lut_1949_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1949_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1949_ff <= lut_1949_out;
            end
        end
        
        assign out_data[1949] = lut_1949_ff;
    end
    else begin : no_ff_1949
        assign out_data[1949] = lut_1949_out;
    end
    endgenerate
    
    
    
    // LUT : 1950
    wire [63:0] lut_1950_table = 64'b0101010101011111010101010101010100000000000000000000000000000000;
    wire [5:0] lut_1950_select = {
                             in_data[401],
                             in_data[614],
                             in_data[61],
                             in_data[764],
                             in_data[45],
                             in_data[151]};
    
    wire lut_1950_out = lut_1950_table[lut_1950_select];
    
    generate
    if ( USE_REG ) begin : ff_1950
        reg   lut_1950_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1950_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1950_ff <= lut_1950_out;
            end
        end
        
        assign out_data[1950] = lut_1950_ff;
    end
    else begin : no_ff_1950
        assign out_data[1950] = lut_1950_out;
    end
    endgenerate
    
    
    
    // LUT : 1951
    wire [63:0] lut_1951_table = 64'b1010101010101010101010101010101011111111111111111111111011111111;
    wire [5:0] lut_1951_select = {
                             in_data[269],
                             in_data[168],
                             in_data[735],
                             in_data[560],
                             in_data[737],
                             in_data[360]};
    
    wire lut_1951_out = lut_1951_table[lut_1951_select];
    
    generate
    if ( USE_REG ) begin : ff_1951
        reg   lut_1951_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1951_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1951_ff <= lut_1951_out;
            end
        end
        
        assign out_data[1951] = lut_1951_ff;
    end
    else begin : no_ff_1951
        assign out_data[1951] = lut_1951_out;
    end
    endgenerate
    
    
    
    // LUT : 1952
    wire [63:0] lut_1952_table = 64'b1111111111111111101010101010101011111111111111110010001000000010;
    wire [5:0] lut_1952_select = {
                             in_data[230],
                             in_data[318],
                             in_data[742],
                             in_data[13],
                             in_data[388],
                             in_data[496]};
    
    wire lut_1952_out = lut_1952_table[lut_1952_select];
    
    generate
    if ( USE_REG ) begin : ff_1952
        reg   lut_1952_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1952_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1952_ff <= lut_1952_out;
            end
        end
        
        assign out_data[1952] = lut_1952_ff;
    end
    else begin : no_ff_1952
        assign out_data[1952] = lut_1952_out;
    end
    endgenerate
    
    
    
    // LUT : 1953
    wire [63:0] lut_1953_table = 64'b0001000100010001000000000000000000010001000100010001000100010001;
    wire [5:0] lut_1953_select = {
                             in_data[355],
                             in_data[383],
                             in_data[703],
                             in_data[309],
                             in_data[687],
                             in_data[630]};
    
    wire lut_1953_out = lut_1953_table[lut_1953_select];
    
    generate
    if ( USE_REG ) begin : ff_1953
        reg   lut_1953_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1953_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1953_ff <= lut_1953_out;
            end
        end
        
        assign out_data[1953] = lut_1953_ff;
    end
    else begin : no_ff_1953
        assign out_data[1953] = lut_1953_out;
    end
    endgenerate
    
    
    
    // LUT : 1954
    wire [63:0] lut_1954_table = 64'b0000000000000000000000000000000000001100000000000000110000001110;
    wire [5:0] lut_1954_select = {
                             in_data[99],
                             in_data[94],
                             in_data[513],
                             in_data[528],
                             in_data[292],
                             in_data[75]};
    
    wire lut_1954_out = lut_1954_table[lut_1954_select];
    
    generate
    if ( USE_REG ) begin : ff_1954
        reg   lut_1954_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1954_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1954_ff <= lut_1954_out;
            end
        end
        
        assign out_data[1954] = lut_1954_ff;
    end
    else begin : no_ff_1954
        assign out_data[1954] = lut_1954_out;
    end
    endgenerate
    
    
    
    // LUT : 1955
    wire [63:0] lut_1955_table = 64'b0000000010110000000000001011000000010000111100010000000011110000;
    wire [5:0] lut_1955_select = {
                             in_data[247],
                             in_data[574],
                             in_data[525],
                             in_data[384],
                             in_data[162],
                             in_data[597]};
    
    wire lut_1955_out = lut_1955_table[lut_1955_select];
    
    generate
    if ( USE_REG ) begin : ff_1955
        reg   lut_1955_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1955_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1955_ff <= lut_1955_out;
            end
        end
        
        assign out_data[1955] = lut_1955_ff;
    end
    else begin : no_ff_1955
        assign out_data[1955] = lut_1955_out;
    end
    endgenerate
    
    
    
    // LUT : 1956
    wire [63:0] lut_1956_table = 64'b0101010101010101010101010101010101110111011101110111011101110111;
    wire [5:0] lut_1956_select = {
                             in_data[494],
                             in_data[84],
                             in_data[198],
                             in_data[765],
                             in_data[542],
                             in_data[488]};
    
    wire lut_1956_out = lut_1956_table[lut_1956_select];
    
    generate
    if ( USE_REG ) begin : ff_1956
        reg   lut_1956_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1956_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1956_ff <= lut_1956_out;
            end
        end
        
        assign out_data[1956] = lut_1956_ff;
    end
    else begin : no_ff_1956
        assign out_data[1956] = lut_1956_out;
    end
    endgenerate
    
    
    
    // LUT : 1957
    wire [63:0] lut_1957_table = 64'b0001010101010111000100010101110100110011101100111001000110111001;
    wire [5:0] lut_1957_select = {
                             in_data[288],
                             in_data[385],
                             in_data[442],
                             in_data[149],
                             in_data[456],
                             in_data[158]};
    
    wire lut_1957_out = lut_1957_table[lut_1957_select];
    
    generate
    if ( USE_REG ) begin : ff_1957
        reg   lut_1957_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1957_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1957_ff <= lut_1957_out;
            end
        end
        
        assign out_data[1957] = lut_1957_ff;
    end
    else begin : no_ff_1957
        assign out_data[1957] = lut_1957_out;
    end
    endgenerate
    
    
    
    // LUT : 1958
    wire [63:0] lut_1958_table = 64'b0000000000000000000000000000000000000000000000000101010101010101;
    wire [5:0] lut_1958_select = {
                             in_data[343],
                             in_data[276],
                             in_data[363],
                             in_data[70],
                             in_data[270],
                             in_data[374]};
    
    wire lut_1958_out = lut_1958_table[lut_1958_select];
    
    generate
    if ( USE_REG ) begin : ff_1958
        reg   lut_1958_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1958_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1958_ff <= lut_1958_out;
            end
        end
        
        assign out_data[1958] = lut_1958_ff;
    end
    else begin : no_ff_1958
        assign out_data[1958] = lut_1958_out;
    end
    endgenerate
    
    
    
    // LUT : 1959
    wire [63:0] lut_1959_table = 64'b1110110011111111110011001100110011111111111111111100110011001100;
    wire [5:0] lut_1959_select = {
                             in_data[390],
                             in_data[426],
                             in_data[46],
                             in_data[224],
                             in_data[423],
                             in_data[167]};
    
    wire lut_1959_out = lut_1959_table[lut_1959_select];
    
    generate
    if ( USE_REG ) begin : ff_1959
        reg   lut_1959_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1959_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1959_ff <= lut_1959_out;
            end
        end
        
        assign out_data[1959] = lut_1959_ff;
    end
    else begin : no_ff_1959
        assign out_data[1959] = lut_1959_out;
    end
    endgenerate
    
    
    
    // LUT : 1960
    wire [63:0] lut_1960_table = 64'b0011001100000000000000000000000000110011001100110000000000000000;
    wire [5:0] lut_1960_select = {
                             in_data[592],
                             in_data[572],
                             in_data[690],
                             in_data[42],
                             in_data[273],
                             in_data[27]};
    
    wire lut_1960_out = lut_1960_table[lut_1960_select];
    
    generate
    if ( USE_REG ) begin : ff_1960
        reg   lut_1960_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1960_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1960_ff <= lut_1960_out;
            end
        end
        
        assign out_data[1960] = lut_1960_ff;
    end
    else begin : no_ff_1960
        assign out_data[1960] = lut_1960_out;
    end
    endgenerate
    
    
    
    // LUT : 1961
    wire [63:0] lut_1961_table = 64'b1111111111111111101110111011101011111111111111111011101110101010;
    wire [5:0] lut_1961_select = {
                             in_data[8],
                             in_data[745],
                             in_data[337],
                             in_data[307],
                             in_data[536],
                             in_data[189]};
    
    wire lut_1961_out = lut_1961_table[lut_1961_select];
    
    generate
    if ( USE_REG ) begin : ff_1961
        reg   lut_1961_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1961_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1961_ff <= lut_1961_out;
            end
        end
        
        assign out_data[1961] = lut_1961_ff;
    end
    else begin : no_ff_1961
        assign out_data[1961] = lut_1961_out;
    end
    endgenerate
    
    
    
    // LUT : 1962
    wire [63:0] lut_1962_table = 64'b0001011100010111001111110111111100000000000000000001000000000000;
    wire [5:0] lut_1962_select = {
                             in_data[348],
                             in_data[263],
                             in_data[68],
                             in_data[605],
                             in_data[340],
                             in_data[321]};
    
    wire lut_1962_out = lut_1962_table[lut_1962_select];
    
    generate
    if ( USE_REG ) begin : ff_1962
        reg   lut_1962_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1962_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1962_ff <= lut_1962_out;
            end
        end
        
        assign out_data[1962] = lut_1962_ff;
    end
    else begin : no_ff_1962
        assign out_data[1962] = lut_1962_out;
    end
    endgenerate
    
    
    
    // LUT : 1963
    wire [63:0] lut_1963_table = 64'b0000101010101010000010101010101010101010101010101010101010101010;
    wire [5:0] lut_1963_select = {
                             in_data[710],
                             in_data[7],
                             in_data[66],
                             in_data[425],
                             in_data[53],
                             in_data[581]};
    
    wire lut_1963_out = lut_1963_table[lut_1963_select];
    
    generate
    if ( USE_REG ) begin : ff_1963
        reg   lut_1963_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1963_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1963_ff <= lut_1963_out;
            end
        end
        
        assign out_data[1963] = lut_1963_ff;
    end
    else begin : no_ff_1963
        assign out_data[1963] = lut_1963_out;
    end
    endgenerate
    
    
    
    // LUT : 1964
    wire [63:0] lut_1964_table = 64'b1111101110111011001000010000001111111011101110110010000100000011;
    wire [5:0] lut_1964_select = {
                             in_data[85],
                             in_data[720],
                             in_data[72],
                             in_data[540],
                             in_data[638],
                             in_data[233]};
    
    wire lut_1964_out = lut_1964_table[lut_1964_select];
    
    generate
    if ( USE_REG ) begin : ff_1964
        reg   lut_1964_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1964_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1964_ff <= lut_1964_out;
            end
        end
        
        assign out_data[1964] = lut_1964_ff;
    end
    else begin : no_ff_1964
        assign out_data[1964] = lut_1964_out;
    end
    endgenerate
    
    
    
    // LUT : 1965
    wire [63:0] lut_1965_table = 64'b0000000000000000101010101010101000000000000000001111111111111111;
    wire [5:0] lut_1965_select = {
                             in_data[668],
                             in_data[602],
                             in_data[734],
                             in_data[83],
                             in_data[335],
                             in_data[316]};
    
    wire lut_1965_out = lut_1965_table[lut_1965_select];
    
    generate
    if ( USE_REG ) begin : ff_1965
        reg   lut_1965_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1965_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1965_ff <= lut_1965_out;
            end
        end
        
        assign out_data[1965] = lut_1965_ff;
    end
    else begin : no_ff_1965
        assign out_data[1965] = lut_1965_out;
    end
    endgenerate
    
    
    
    // LUT : 1966
    wire [63:0] lut_1966_table = 64'b1011101000000000101110100000000011111111100110011111111111111111;
    wire [5:0] lut_1966_select = {
                             in_data[290],
                             in_data[274],
                             in_data[651],
                             in_data[391],
                             in_data[470],
                             in_data[544]};
    
    wire lut_1966_out = lut_1966_table[lut_1966_select];
    
    generate
    if ( USE_REG ) begin : ff_1966
        reg   lut_1966_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1966_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1966_ff <= lut_1966_out;
            end
        end
        
        assign out_data[1966] = lut_1966_ff;
    end
    else begin : no_ff_1966
        assign out_data[1966] = lut_1966_out;
    end
    endgenerate
    
    
    
    // LUT : 1967
    wire [63:0] lut_1967_table = 64'b0000000011110000000000001111000000000000111100000000000011110000;
    wire [5:0] lut_1967_select = {
                             in_data[700],
                             in_data[82],
                             in_data[125],
                             in_data[326],
                             in_data[109],
                             in_data[107]};
    
    wire lut_1967_out = lut_1967_table[lut_1967_select];
    
    generate
    if ( USE_REG ) begin : ff_1967
        reg   lut_1967_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1967_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1967_ff <= lut_1967_out;
            end
        end
        
        assign out_data[1967] = lut_1967_ff;
    end
    else begin : no_ff_1967
        assign out_data[1967] = lut_1967_out;
    end
    endgenerate
    
    
    
    // LUT : 1968
    wire [63:0] lut_1968_table = 64'b1111000011110000010111000101110110111110101110110000100000001010;
    wire [5:0] lut_1968_select = {
                             in_data[431],
                             in_data[406],
                             in_data[248],
                             in_data[486],
                             in_data[666],
                             in_data[520]};
    
    wire lut_1968_out = lut_1968_table[lut_1968_select];
    
    generate
    if ( USE_REG ) begin : ff_1968
        reg   lut_1968_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1968_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1968_ff <= lut_1968_out;
            end
        end
        
        assign out_data[1968] = lut_1968_ff;
    end
    else begin : no_ff_1968
        assign out_data[1968] = lut_1968_out;
    end
    endgenerate
    
    
    
    // LUT : 1969
    wire [63:0] lut_1969_table = 64'b1111111111111111111111111111111111001110110011111111110011001100;
    wire [5:0] lut_1969_select = {
                             in_data[325],
                             in_data[150],
                             in_data[633],
                             in_data[371],
                             in_data[103],
                             in_data[759]};
    
    wire lut_1969_out = lut_1969_table[lut_1969_select];
    
    generate
    if ( USE_REG ) begin : ff_1969
        reg   lut_1969_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1969_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1969_ff <= lut_1969_out;
            end
        end
        
        assign out_data[1969] = lut_1969_ff;
    end
    else begin : no_ff_1969
        assign out_data[1969] = lut_1969_out;
    end
    endgenerate
    
    
    
    // LUT : 1970
    wire [63:0] lut_1970_table = 64'b1100000000000101111000100010001111000111000001111110111100000011;
    wire [5:0] lut_1970_select = {
                             in_data[291],
                             in_data[132],
                             in_data[234],
                             in_data[370],
                             in_data[482],
                             in_data[328]};
    
    wire lut_1970_out = lut_1970_table[lut_1970_select];
    
    generate
    if ( USE_REG ) begin : ff_1970
        reg   lut_1970_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1970_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1970_ff <= lut_1970_out;
            end
        end
        
        assign out_data[1970] = lut_1970_ff;
    end
    else begin : no_ff_1970
        assign out_data[1970] = lut_1970_out;
    end
    endgenerate
    
    
    
    // LUT : 1971
    wire [63:0] lut_1971_table = 64'b0000000000000000111111111100000011111111111111111111111111111111;
    wire [5:0] lut_1971_select = {
                             in_data[429],
                             in_data[331],
                             in_data[539],
                             in_data[361],
                             in_data[40],
                             in_data[449]};
    
    wire lut_1971_out = lut_1971_table[lut_1971_select];
    
    generate
    if ( USE_REG ) begin : ff_1971
        reg   lut_1971_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1971_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1971_ff <= lut_1971_out;
            end
        end
        
        assign out_data[1971] = lut_1971_ff;
    end
    else begin : no_ff_1971
        assign out_data[1971] = lut_1971_out;
    end
    endgenerate
    
    
    
    // LUT : 1972
    wire [63:0] lut_1972_table = 64'b1101110100000000110111010000000011111111110101011111111111011101;
    wire [5:0] lut_1972_select = {
                             in_data[517],
                             in_data[559],
                             in_data[372],
                             in_data[48],
                             in_data[506],
                             in_data[601]};
    
    wire lut_1972_out = lut_1972_table[lut_1972_select];
    
    generate
    if ( USE_REG ) begin : ff_1972
        reg   lut_1972_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1972_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1972_ff <= lut_1972_out;
            end
        end
        
        assign out_data[1972] = lut_1972_ff;
    end
    else begin : no_ff_1972
        assign out_data[1972] = lut_1972_out;
    end
    endgenerate
    
    
    
    // LUT : 1973
    wire [63:0] lut_1973_table = 64'b0000000000000000000000000000000010101010101110111010001010111011;
    wire [5:0] lut_1973_select = {
                             in_data[686],
                             in_data[10],
                             in_data[159],
                             in_data[188],
                             in_data[283],
                             in_data[747]};
    
    wire lut_1973_out = lut_1973_table[lut_1973_select];
    
    generate
    if ( USE_REG ) begin : ff_1973
        reg   lut_1973_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1973_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1973_ff <= lut_1973_out;
            end
        end
        
        assign out_data[1973] = lut_1973_ff;
    end
    else begin : no_ff_1973
        assign out_data[1973] = lut_1973_out;
    end
    endgenerate
    
    
    
    // LUT : 1974
    wire [63:0] lut_1974_table = 64'b0000000010111010111111111111111100000000000000001111010111110000;
    wire [5:0] lut_1974_select = {
                             in_data[246],
                             in_data[610],
                             in_data[603],
                             in_data[203],
                             in_data[751],
                             in_data[262]};
    
    wire lut_1974_out = lut_1974_table[lut_1974_select];
    
    generate
    if ( USE_REG ) begin : ff_1974
        reg   lut_1974_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1974_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1974_ff <= lut_1974_out;
            end
        end
        
        assign out_data[1974] = lut_1974_ff;
    end
    else begin : no_ff_1974
        assign out_data[1974] = lut_1974_out;
    end
    endgenerate
    
    
    
    // LUT : 1975
    wire [63:0] lut_1975_table = 64'b0000011100000111000000010000000100000111000011110000001100000011;
    wire [5:0] lut_1975_select = {
                             in_data[718],
                             in_data[367],
                             in_data[615],
                             in_data[659],
                             in_data[537],
                             in_data[691]};
    
    wire lut_1975_out = lut_1975_table[lut_1975_select];
    
    generate
    if ( USE_REG ) begin : ff_1975
        reg   lut_1975_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1975_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1975_ff <= lut_1975_out;
            end
        end
        
        assign out_data[1975] = lut_1975_ff;
    end
    else begin : no_ff_1975
        assign out_data[1975] = lut_1975_out;
    end
    endgenerate
    
    
    
    // LUT : 1976
    wire [63:0] lut_1976_table = 64'b0000000000000000000100010000000000110011000000000011001100110011;
    wire [5:0] lut_1976_select = {
                             in_data[556],
                             in_data[467],
                             in_data[621],
                             in_data[476],
                             in_data[95],
                             in_data[761]};
    
    wire lut_1976_out = lut_1976_table[lut_1976_select];
    
    generate
    if ( USE_REG ) begin : ff_1976
        reg   lut_1976_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1976_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1976_ff <= lut_1976_out;
            end
        end
        
        assign out_data[1976] = lut_1976_ff;
    end
    else begin : no_ff_1976
        assign out_data[1976] = lut_1976_out;
    end
    endgenerate
    
    
    
    // LUT : 1977
    wire [63:0] lut_1977_table = 64'b1011111110101111101111111011111110101111101011111010111110101111;
    wire [5:0] lut_1977_select = {
                             in_data[108],
                             in_data[16],
                             in_data[669],
                             in_data[485],
                             in_data[588],
                             in_data[164]};
    
    wire lut_1977_out = lut_1977_table[lut_1977_select];
    
    generate
    if ( USE_REG ) begin : ff_1977
        reg   lut_1977_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1977_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1977_ff <= lut_1977_out;
            end
        end
        
        assign out_data[1977] = lut_1977_ff;
    end
    else begin : no_ff_1977
        assign out_data[1977] = lut_1977_out;
    end
    endgenerate
    
    
    
    // LUT : 1978
    wire [63:0] lut_1978_table = 64'b1100110011001100110011001100110011001100110111001110100011001100;
    wire [5:0] lut_1978_select = {
                             in_data[0],
                             in_data[129],
                             in_data[301],
                             in_data[421],
                             in_data[214],
                             in_data[235]};
    
    wire lut_1978_out = lut_1978_table[lut_1978_select];
    
    generate
    if ( USE_REG ) begin : ff_1978
        reg   lut_1978_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1978_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1978_ff <= lut_1978_out;
            end
        end
        
        assign out_data[1978] = lut_1978_ff;
    end
    else begin : no_ff_1978
        assign out_data[1978] = lut_1978_out;
    end
    endgenerate
    
    
    
    // LUT : 1979
    wire [63:0] lut_1979_table = 64'b1111111111001100110011000000000011111111111111111111111111001100;
    wire [5:0] lut_1979_select = {
                             in_data[220],
                             in_data[411],
                             in_data[257],
                             in_data[166],
                             in_data[611],
                             in_data[339]};
    
    wire lut_1979_out = lut_1979_table[lut_1979_select];
    
    generate
    if ( USE_REG ) begin : ff_1979
        reg   lut_1979_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1979_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1979_ff <= lut_1979_out;
            end
        end
        
        assign out_data[1979] = lut_1979_ff;
    end
    else begin : no_ff_1979
        assign out_data[1979] = lut_1979_out;
    end
    endgenerate
    
    
    
    // LUT : 1980
    wire [63:0] lut_1980_table = 64'b1111111111110001111111110101000011111111111101011111111101010000;
    wire [5:0] lut_1980_select = {
                             in_data[113],
                             in_data[445],
                             in_data[595],
                             in_data[239],
                             in_data[240],
                             in_data[693]};
    
    wire lut_1980_out = lut_1980_table[lut_1980_select];
    
    generate
    if ( USE_REG ) begin : ff_1980
        reg   lut_1980_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1980_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1980_ff <= lut_1980_out;
            end
        end
        
        assign out_data[1980] = lut_1980_ff;
    end
    else begin : no_ff_1980
        assign out_data[1980] = lut_1980_out;
    end
    endgenerate
    
    
    
    // LUT : 1981
    wire [63:0] lut_1981_table = 64'b0011001100100011101110111010101100110011001000110010101100100010;
    wire [5:0] lut_1981_select = {
                             in_data[632],
                             in_data[608],
                             in_data[530],
                             in_data[714],
                             in_data[342],
                             in_data[71]};
    
    wire lut_1981_out = lut_1981_table[lut_1981_select];
    
    generate
    if ( USE_REG ) begin : ff_1981
        reg   lut_1981_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1981_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1981_ff <= lut_1981_out;
            end
        end
        
        assign out_data[1981] = lut_1981_ff;
    end
    else begin : no_ff_1981
        assign out_data[1981] = lut_1981_out;
    end
    endgenerate
    
    
    
    // LUT : 1982
    wire [63:0] lut_1982_table = 64'b0101010100000000010101010100010011010101000000001111111101000100;
    wire [5:0] lut_1982_select = {
                             in_data[504],
                             in_data[620],
                             in_data[683],
                             in_data[475],
                             in_data[619],
                             in_data[131]};
    
    wire lut_1982_out = lut_1982_table[lut_1982_select];
    
    generate
    if ( USE_REG ) begin : ff_1982
        reg   lut_1982_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1982_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1982_ff <= lut_1982_out;
            end
        end
        
        assign out_data[1982] = lut_1982_ff;
    end
    else begin : no_ff_1982
        assign out_data[1982] = lut_1982_out;
    end
    endgenerate
    
    
    
    // LUT : 1983
    wire [63:0] lut_1983_table = 64'b0000000000000000001100110011001100110011001100110011001100110011;
    wire [5:0] lut_1983_select = {
                             in_data[354],
                             in_data[294],
                             in_data[59],
                             in_data[365],
                             in_data[241],
                             in_data[139]};
    
    wire lut_1983_out = lut_1983_table[lut_1983_select];
    
    generate
    if ( USE_REG ) begin : ff_1983
        reg   lut_1983_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1983_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1983_ff <= lut_1983_out;
            end
        end
        
        assign out_data[1983] = lut_1983_ff;
    end
    else begin : no_ff_1983
        assign out_data[1983] = lut_1983_out;
    end
    endgenerate
    
    
    
    // LUT : 1984
    wire [63:0] lut_1984_table = 64'b1111111111111111111111110000000011111111111011111111111100000000;
    wire [5:0] lut_1984_select = {
                             in_data[112],
                             in_data[571],
                             in_data[529],
                             in_data[101],
                             in_data[422],
                             in_data[725]};
    
    wire lut_1984_out = lut_1984_table[lut_1984_select];
    
    generate
    if ( USE_REG ) begin : ff_1984
        reg   lut_1984_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1984_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1984_ff <= lut_1984_out;
            end
        end
        
        assign out_data[1984] = lut_1984_ff;
    end
    else begin : no_ff_1984
        assign out_data[1984] = lut_1984_out;
    end
    endgenerate
    
    
    
    // LUT : 1985
    wire [63:0] lut_1985_table = 64'b1100010100000100111111111100110111000101000000001111111111001101;
    wire [5:0] lut_1985_select = {
                             in_data[138],
                             in_data[192],
                             in_data[39],
                             in_data[437],
                             in_data[64],
                             in_data[705]};
    
    wire lut_1985_out = lut_1985_table[lut_1985_select];
    
    generate
    if ( USE_REG ) begin : ff_1985
        reg   lut_1985_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1985_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1985_ff <= lut_1985_out;
            end
        end
        
        assign out_data[1985] = lut_1985_ff;
    end
    else begin : no_ff_1985
        assign out_data[1985] = lut_1985_out;
    end
    endgenerate
    
    
    
    // LUT : 1986
    wire [63:0] lut_1986_table = 64'b0000000001001101000000000100110100000000010011010000000011001101;
    wire [5:0] lut_1986_select = {
                             in_data[51],
                             in_data[769],
                             in_data[204],
                             in_data[92],
                             in_data[277],
                             in_data[207]};
    
    wire lut_1986_out = lut_1986_table[lut_1986_select];
    
    generate
    if ( USE_REG ) begin : ff_1986
        reg   lut_1986_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1986_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1986_ff <= lut_1986_out;
            end
        end
        
        assign out_data[1986] = lut_1986_ff;
    end
    else begin : no_ff_1986
        assign out_data[1986] = lut_1986_out;
    end
    endgenerate
    
    
    
    // LUT : 1987
    wire [63:0] lut_1987_table = 64'b1111111111111111011100011111111100000000111111110000000011111111;
    wire [5:0] lut_1987_select = {
                             in_data[208],
                             in_data[667],
                             in_data[323],
                             in_data[733],
                             in_data[473],
                             in_data[261]};
    
    wire lut_1987_out = lut_1987_table[lut_1987_select];
    
    generate
    if ( USE_REG ) begin : ff_1987
        reg   lut_1987_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1987_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1987_ff <= lut_1987_out;
            end
        end
        
        assign out_data[1987] = lut_1987_ff;
    end
    else begin : no_ff_1987
        assign out_data[1987] = lut_1987_out;
    end
    endgenerate
    
    
    
    // LUT : 1988
    wire [63:0] lut_1988_table = 64'b1111001111111111111100111111111100110000001100000011000000110010;
    wire [5:0] lut_1988_select = {
                             in_data[229],
                             in_data[250],
                             in_data[359],
                             in_data[661],
                             in_data[299],
                             in_data[9]};
    
    wire lut_1988_out = lut_1988_table[lut_1988_select];
    
    generate
    if ( USE_REG ) begin : ff_1988
        reg   lut_1988_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1988_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1988_ff <= lut_1988_out;
            end
        end
        
        assign out_data[1988] = lut_1988_ff;
    end
    else begin : no_ff_1988
        assign out_data[1988] = lut_1988_out;
    end
    endgenerate
    
    
    
    // LUT : 1989
    wire [63:0] lut_1989_table = 64'b1110111010001000111111111100111111101111100010101111111111101111;
    wire [5:0] lut_1989_select = {
                             in_data[54],
                             in_data[97],
                             in_data[171],
                             in_data[706],
                             in_data[450],
                             in_data[642]};
    
    wire lut_1989_out = lut_1989_table[lut_1989_select];
    
    generate
    if ( USE_REG ) begin : ff_1989
        reg   lut_1989_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1989_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1989_ff <= lut_1989_out;
            end
        end
        
        assign out_data[1989] = lut_1989_ff;
    end
    else begin : no_ff_1989
        assign out_data[1989] = lut_1989_out;
    end
    endgenerate
    
    
    
    // LUT : 1990
    wire [63:0] lut_1990_table = 64'b1111001111110010111100111111001100110000001100001011000010110001;
    wire [5:0] lut_1990_select = {
                             in_data[440],
                             in_data[78],
                             in_data[746],
                             in_data[567],
                             in_data[128],
                             in_data[134]};
    
    wire lut_1990_out = lut_1990_table[lut_1990_select];
    
    generate
    if ( USE_REG ) begin : ff_1990
        reg   lut_1990_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1990_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1990_ff <= lut_1990_out;
            end
        end
        
        assign out_data[1990] = lut_1990_ff;
    end
    else begin : no_ff_1990
        assign out_data[1990] = lut_1990_out;
    end
    endgenerate
    
    
    
    // LUT : 1991
    wire [63:0] lut_1991_table = 64'b0000000000000000100000100000000000000000000000001010101110101011;
    wire [5:0] lut_1991_select = {
                             in_data[443],
                             in_data[286],
                             in_data[753],
                             in_data[748],
                             in_data[489],
                             in_data[490]};
    
    wire lut_1991_out = lut_1991_table[lut_1991_select];
    
    generate
    if ( USE_REG ) begin : ff_1991
        reg   lut_1991_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1991_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1991_ff <= lut_1991_out;
            end
        end
        
        assign out_data[1991] = lut_1991_ff;
    end
    else begin : no_ff_1991
        assign out_data[1991] = lut_1991_out;
    end
    endgenerate
    
    
    
    // LUT : 1992
    wire [63:0] lut_1992_table = 64'b1111111111111111110011100000110011111111111111111100111000001100;
    wire [5:0] lut_1992_select = {
                             in_data[676],
                             in_data[433],
                             in_data[598],
                             in_data[427],
                             in_data[120],
                             in_data[38]};
    
    wire lut_1992_out = lut_1992_table[lut_1992_select];
    
    generate
    if ( USE_REG ) begin : ff_1992
        reg   lut_1992_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1992_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1992_ff <= lut_1992_out;
            end
        end
        
        assign out_data[1992] = lut_1992_ff;
    end
    else begin : no_ff_1992
        assign out_data[1992] = lut_1992_out;
    end
    endgenerate
    
    
    
    // LUT : 1993
    wire [63:0] lut_1993_table = 64'b1100110011011100110011001100110011001100110011001100110011001100;
    wire [5:0] lut_1993_select = {
                             in_data[80],
                             in_data[557],
                             in_data[18],
                             in_data[664],
                             in_data[213],
                             in_data[709]};
    
    wire lut_1993_out = lut_1993_table[lut_1993_select];
    
    generate
    if ( USE_REG ) begin : ff_1993
        reg   lut_1993_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1993_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1993_ff <= lut_1993_out;
            end
        end
        
        assign out_data[1993] = lut_1993_ff;
    end
    else begin : no_ff_1993
        assign out_data[1993] = lut_1993_out;
    end
    endgenerate
    
    
    
    // LUT : 1994
    wire [63:0] lut_1994_table = 64'b0001000100010001000000000001000100010001000100010000000000010001;
    wire [5:0] lut_1994_select = {
                             in_data[701],
                             in_data[12],
                             in_data[732],
                             in_data[23],
                             in_data[623],
                             in_data[749]};
    
    wire lut_1994_out = lut_1994_table[lut_1994_select];
    
    generate
    if ( USE_REG ) begin : ff_1994
        reg   lut_1994_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1994_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1994_ff <= lut_1994_out;
            end
        end
        
        assign out_data[1994] = lut_1994_ff;
    end
    else begin : no_ff_1994
        assign out_data[1994] = lut_1994_out;
    end
    endgenerate
    
    
    
    // LUT : 1995
    wire [63:0] lut_1995_table = 64'b0000000000000000000000000000000000000000000000000001000100010001;
    wire [5:0] lut_1995_select = {
                             in_data[527],
                             in_data[554],
                             in_data[546],
                             in_data[757],
                             in_data[452],
                             in_data[152]};
    
    wire lut_1995_out = lut_1995_table[lut_1995_select];
    
    generate
    if ( USE_REG ) begin : ff_1995
        reg   lut_1995_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1995_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1995_ff <= lut_1995_out;
            end
        end
        
        assign out_data[1995] = lut_1995_ff;
    end
    else begin : no_ff_1995
        assign out_data[1995] = lut_1995_out;
    end
    endgenerate
    
    
    
    // LUT : 1996
    wire [63:0] lut_1996_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_1996_select = {
                             in_data[57],
                             in_data[211],
                             in_data[781],
                             in_data[119],
                             in_data[34],
                             in_data[377]};
    
    wire lut_1996_out = lut_1996_table[lut_1996_select];
    
    generate
    if ( USE_REG ) begin : ff_1996
        reg   lut_1996_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1996_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1996_ff <= lut_1996_out;
            end
        end
        
        assign out_data[1996] = lut_1996_ff;
    end
    else begin : no_ff_1996
        assign out_data[1996] = lut_1996_out;
    end
    endgenerate
    
    
    
    // LUT : 1997
    wire [63:0] lut_1997_table = 64'b0100000000000000010000000000000011111111110111001111111111010101;
    wire [5:0] lut_1997_select = {
                             in_data[330],
                             in_data[266],
                             in_data[160],
                             in_data[105],
                             in_data[639],
                             in_data[314]};
    
    wire lut_1997_out = lut_1997_table[lut_1997_select];
    
    generate
    if ( USE_REG ) begin : ff_1997
        reg   lut_1997_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1997_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1997_ff <= lut_1997_out;
            end
        end
        
        assign out_data[1997] = lut_1997_ff;
    end
    else begin : no_ff_1997
        assign out_data[1997] = lut_1997_out;
    end
    endgenerate
    
    
    
    // LUT : 1998
    wire [63:0] lut_1998_table = 64'b0111011101110111111111110111011111111111011111111111111100000000;
    wire [5:0] lut_1998_select = {
                             in_data[606],
                             in_data[553],
                             in_data[416],
                             in_data[22],
                             in_data[479],
                             in_data[175]};
    
    wire lut_1998_out = lut_1998_table[lut_1998_select];
    
    generate
    if ( USE_REG ) begin : ff_1998
        reg   lut_1998_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1998_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1998_ff <= lut_1998_out;
            end
        end
        
        assign out_data[1998] = lut_1998_ff;
    end
    else begin : no_ff_1998
        assign out_data[1998] = lut_1998_out;
    end
    endgenerate
    
    
    
    // LUT : 1999
    wire [63:0] lut_1999_table = 64'b0000000000000000000000000000000011111111111111111111111100110011;
    wire [5:0] lut_1999_select = {
                             in_data[387],
                             in_data[311],
                             in_data[313],
                             in_data[503],
                             in_data[591],
                             in_data[55]};
    
    wire lut_1999_out = lut_1999_table[lut_1999_select];
    
    generate
    if ( USE_REG ) begin : ff_1999
        reg   lut_1999_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1999_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1999_ff <= lut_1999_out;
            end
        end
        
        assign out_data[1999] = lut_1999_ff;
    end
    else begin : no_ff_1999
        assign out_data[1999] = lut_1999_out;
    end
    endgenerate
    
    
    
    // LUT : 2000
    wire [63:0] lut_2000_table = 64'b0000110100001101010011010100110100001101000011010100110101001101;
    wire [5:0] lut_2000_select = {
                             in_data[739],
                             in_data[565],
                             in_data[675],
                             in_data[153],
                             in_data[217],
                             in_data[76]};
    
    wire lut_2000_out = lut_2000_table[lut_2000_select];
    
    generate
    if ( USE_REG ) begin : ff_2000
        reg   lut_2000_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2000_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2000_ff <= lut_2000_out;
            end
        end
        
        assign out_data[2000] = lut_2000_ff;
    end
    else begin : no_ff_2000
        assign out_data[2000] = lut_2000_out;
    end
    endgenerate
    
    
    
    // LUT : 2001
    wire [63:0] lut_2001_table = 64'b0101110111010101111111111111111101010101010101010101010101010101;
    wire [5:0] lut_2001_select = {
                             in_data[260],
                             in_data[770],
                             in_data[310],
                             in_data[28],
                             in_data[695],
                             in_data[350]};
    
    wire lut_2001_out = lut_2001_table[lut_2001_select];
    
    generate
    if ( USE_REG ) begin : ff_2001
        reg   lut_2001_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2001_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2001_ff <= lut_2001_out;
            end
        end
        
        assign out_data[2001] = lut_2001_ff;
    end
    else begin : no_ff_2001
        assign out_data[2001] = lut_2001_out;
    end
    endgenerate
    
    
    
    // LUT : 2002
    wire [63:0] lut_2002_table = 64'b1111110111111101111111001111110011111111111111111111111111111111;
    wire [5:0] lut_2002_select = {
                             in_data[156],
                             in_data[201],
                             in_data[24],
                             in_data[285],
                             in_data[136],
                             in_data[215]};
    
    wire lut_2002_out = lut_2002_table[lut_2002_select];
    
    generate
    if ( USE_REG ) begin : ff_2002
        reg   lut_2002_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2002_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2002_ff <= lut_2002_out;
            end
        end
        
        assign out_data[2002] = lut_2002_ff;
    end
    else begin : no_ff_2002
        assign out_data[2002] = lut_2002_out;
    end
    endgenerate
    
    
    
    // LUT : 2003
    wire [63:0] lut_2003_table = 64'b1111000011111000000000001111000011110000111110000000000011110000;
    wire [5:0] lut_2003_select = {
                             in_data[32],
                             in_data[243],
                             in_data[127],
                             in_data[628],
                             in_data[727],
                             in_data[147]};
    
    wire lut_2003_out = lut_2003_table[lut_2003_select];
    
    generate
    if ( USE_REG ) begin : ff_2003
        reg   lut_2003_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2003_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2003_ff <= lut_2003_out;
            end
        end
        
        assign out_data[2003] = lut_2003_ff;
    end
    else begin : no_ff_2003
        assign out_data[2003] = lut_2003_out;
    end
    endgenerate
    
    
    
    // LUT : 2004
    wire [63:0] lut_2004_table = 64'b1111111111111111111011101110111011111111111111101110111011101110;
    wire [5:0] lut_2004_select = {
                             in_data[62],
                             in_data[122],
                             in_data[766],
                             in_data[523],
                             in_data[100],
                             in_data[516]};
    
    wire lut_2004_out = lut_2004_table[lut_2004_select];
    
    generate
    if ( USE_REG ) begin : ff_2004
        reg   lut_2004_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2004_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2004_ff <= lut_2004_out;
            end
        end
        
        assign out_data[2004] = lut_2004_ff;
    end
    else begin : no_ff_2004
        assign out_data[2004] = lut_2004_out;
    end
    endgenerate
    
    
    
    // LUT : 2005
    wire [63:0] lut_2005_table = 64'b1111001111110011001000110010001111110011101100110010001000100011;
    wire [5:0] lut_2005_select = {
                             in_data[451],
                             in_data[123],
                             in_data[731],
                             in_data[145],
                             in_data[663],
                             in_data[221]};
    
    wire lut_2005_out = lut_2005_table[lut_2005_select];
    
    generate
    if ( USE_REG ) begin : ff_2005
        reg   lut_2005_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2005_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2005_ff <= lut_2005_out;
            end
        end
        
        assign out_data[2005] = lut_2005_ff;
    end
    else begin : no_ff_2005
        assign out_data[2005] = lut_2005_out;
    end
    endgenerate
    
    
    
    // LUT : 2006
    wire [63:0] lut_2006_table = 64'b1111011111111111000100010011001111111111111111110000001100110011;
    wire [5:0] lut_2006_select = {
                             in_data[141],
                             in_data[585],
                             in_data[418],
                             in_data[338],
                             in_data[324],
                             in_data[280]};
    
    wire lut_2006_out = lut_2006_table[lut_2006_select];
    
    generate
    if ( USE_REG ) begin : ff_2006
        reg   lut_2006_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2006_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2006_ff <= lut_2006_out;
            end
        end
        
        assign out_data[2006] = lut_2006_ff;
    end
    else begin : no_ff_2006
        assign out_data[2006] = lut_2006_out;
    end
    endgenerate
    
    
    
    // LUT : 2007
    wire [63:0] lut_2007_table = 64'b1111100111011101111110011101100111011001110101011111100111011001;
    wire [5:0] lut_2007_select = {
                             in_data[341],
                             in_data[96],
                             in_data[511],
                             in_data[332],
                             in_data[272],
                             in_data[322]};
    
    wire lut_2007_out = lut_2007_table[lut_2007_select];
    
    generate
    if ( USE_REG ) begin : ff_2007
        reg   lut_2007_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2007_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2007_ff <= lut_2007_out;
            end
        end
        
        assign out_data[2007] = lut_2007_ff;
    end
    else begin : no_ff_2007
        assign out_data[2007] = lut_2007_out;
    end
    endgenerate
    
    
    
    // LUT : 2008
    wire [63:0] lut_2008_table = 64'b1111111111111111111111111111111111111010111111101111101011111110;
    wire [5:0] lut_2008_select = {
                             in_data[555],
                             in_data[308],
                             in_data[778],
                             in_data[362],
                             in_data[1],
                             in_data[613]};
    
    wire lut_2008_out = lut_2008_table[lut_2008_select];
    
    generate
    if ( USE_REG ) begin : ff_2008
        reg   lut_2008_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2008_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2008_ff <= lut_2008_out;
            end
        end
        
        assign out_data[2008] = lut_2008_ff;
    end
    else begin : no_ff_2008
        assign out_data[2008] = lut_2008_out;
    end
    endgenerate
    
    
    
    // LUT : 2009
    wire [63:0] lut_2009_table = 64'b1111111111110000111111111111010011111111111100001111111111110000;
    wire [5:0] lut_2009_select = {
                             in_data[89],
                             in_data[631],
                             in_data[124],
                             in_data[174],
                             in_data[558],
                             in_data[699]};
    
    wire lut_2009_out = lut_2009_table[lut_2009_select];
    
    generate
    if ( USE_REG ) begin : ff_2009
        reg   lut_2009_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2009_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2009_ff <= lut_2009_out;
            end
        end
        
        assign out_data[2009] = lut_2009_ff;
    end
    else begin : no_ff_2009
        assign out_data[2009] = lut_2009_out;
    end
    endgenerate
    
    
    
    // LUT : 2010
    wire [63:0] lut_2010_table = 64'b0000000000000000000100000101000001010101010101010101010101010101;
    wire [5:0] lut_2010_select = {
                             in_data[509],
                             in_data[643],
                             in_data[783],
                             in_data[656],
                             in_data[29],
                             in_data[434]};
    
    wire lut_2010_out = lut_2010_table[lut_2010_select];
    
    generate
    if ( USE_REG ) begin : ff_2010
        reg   lut_2010_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2010_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2010_ff <= lut_2010_out;
            end
        end
        
        assign out_data[2010] = lut_2010_ff;
    end
    else begin : no_ff_2010
        assign out_data[2010] = lut_2010_out;
    end
    endgenerate
    
    
    
    // LUT : 2011
    wire [63:0] lut_2011_table = 64'b0000001000000010000000000000001100000000000000000011001100110011;
    wire [5:0] lut_2011_select = {
                             in_data[347],
                             in_data[551],
                             in_data[779],
                             in_data[65],
                             in_data[344],
                             in_data[287]};
    
    wire lut_2011_out = lut_2011_table[lut_2011_select];
    
    generate
    if ( USE_REG ) begin : ff_2011
        reg   lut_2011_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2011_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2011_ff <= lut_2011_out;
            end
        end
        
        assign out_data[2011] = lut_2011_ff;
    end
    else begin : no_ff_2011
        assign out_data[2011] = lut_2011_out;
    end
    endgenerate
    
    
    
    // LUT : 2012
    wire [63:0] lut_2012_table = 64'b1100111111001100111011111100110011001111110011001100111111001111;
    wire [5:0] lut_2012_select = {
                             in_data[465],
                             in_data[646],
                             in_data[743],
                             in_data[178],
                             in_data[464],
                             in_data[47]};
    
    wire lut_2012_out = lut_2012_table[lut_2012_select];
    
    generate
    if ( USE_REG ) begin : ff_2012
        reg   lut_2012_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2012_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2012_ff <= lut_2012_out;
            end
        end
        
        assign out_data[2012] = lut_2012_ff;
    end
    else begin : no_ff_2012
        assign out_data[2012] = lut_2012_out;
    end
    endgenerate
    
    
    
    // LUT : 2013
    wire [63:0] lut_2013_table = 64'b1111111111111111111111111111111111111111101010101111111110100010;
    wire [5:0] lut_2013_select = {
                             in_data[104],
                             in_data[730],
                             in_data[255],
                             in_data[21],
                             in_data[74],
                             in_data[413]};
    
    wire lut_2013_out = lut_2013_table[lut_2013_select];
    
    generate
    if ( USE_REG ) begin : ff_2013
        reg   lut_2013_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2013_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2013_ff <= lut_2013_out;
            end
        end
        
        assign out_data[2013] = lut_2013_ff;
    end
    else begin : no_ff_2013
        assign out_data[2013] = lut_2013_out;
    end
    endgenerate
    
    
    
    // LUT : 2014
    wire [63:0] lut_2014_table = 64'b0000000001010100100000001111010111111010111111111010101011111111;
    wire [5:0] lut_2014_select = {
                             in_data[410],
                             in_data[190],
                             in_data[462],
                             in_data[640],
                             in_data[117],
                             in_data[289]};
    
    wire lut_2014_out = lut_2014_table[lut_2014_select];
    
    generate
    if ( USE_REG ) begin : ff_2014
        reg   lut_2014_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2014_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2014_ff <= lut_2014_out;
            end
        end
        
        assign out_data[2014] = lut_2014_ff;
    end
    else begin : no_ff_2014
        assign out_data[2014] = lut_2014_out;
    end
    endgenerate
    
    
    
    // LUT : 2015
    wire [63:0] lut_2015_table = 64'b1111111100001100111111110000110011111111000011001111111100001100;
    wire [5:0] lut_2015_select = {
                             in_data[767],
                             in_data[6],
                             in_data[259],
                             in_data[500],
                             in_data[379],
                             in_data[447]};
    
    wire lut_2015_out = lut_2015_table[lut_2015_select];
    
    generate
    if ( USE_REG ) begin : ff_2015
        reg   lut_2015_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2015_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2015_ff <= lut_2015_out;
            end
        end
        
        assign out_data[2015] = lut_2015_ff;
    end
    else begin : no_ff_2015
        assign out_data[2015] = lut_2015_out;
    end
    endgenerate
    
    
    
    // LUT : 2016
    wire [63:0] lut_2016_table = 64'b0011001100110011000000000000000000010011001100110000000000100000;
    wire [5:0] lut_2016_select = {
                             in_data[704],
                             in_data[300],
                             in_data[146],
                             in_data[172],
                             in_data[405],
                             in_data[90]};
    
    wire lut_2016_out = lut_2016_table[lut_2016_select];
    
    generate
    if ( USE_REG ) begin : ff_2016
        reg   lut_2016_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2016_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2016_ff <= lut_2016_out;
            end
        end
        
        assign out_data[2016] = lut_2016_ff;
    end
    else begin : no_ff_2016
        assign out_data[2016] = lut_2016_out;
    end
    endgenerate
    
    
    
    // LUT : 2017
    wire [63:0] lut_2017_table = 64'b0000111111001111000011111101111100000000110011000000110011001100;
    wire [5:0] lut_2017_select = {
                             in_data[507],
                             in_data[33],
                             in_data[232],
                             in_data[568],
                             in_data[495],
                             in_data[50]};
    
    wire lut_2017_out = lut_2017_table[lut_2017_select];
    
    generate
    if ( USE_REG ) begin : ff_2017
        reg   lut_2017_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2017_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2017_ff <= lut_2017_out;
            end
        end
        
        assign out_data[2017] = lut_2017_ff;
    end
    else begin : no_ff_2017
        assign out_data[2017] = lut_2017_out;
    end
    endgenerate
    
    
    
    // LUT : 2018
    wire [63:0] lut_2018_table = 64'b0000000000000000000000000000000000001111000011110000000000000000;
    wire [5:0] lut_2018_select = {
                             in_data[637],
                             in_data[352],
                             in_data[5],
                             in_data[474],
                             in_data[364],
                             in_data[173]};
    
    wire lut_2018_out = lut_2018_table[lut_2018_select];
    
    generate
    if ( USE_REG ) begin : ff_2018
        reg   lut_2018_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2018_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2018_ff <= lut_2018_out;
            end
        end
        
        assign out_data[2018] = lut_2018_ff;
    end
    else begin : no_ff_2018
        assign out_data[2018] = lut_2018_out;
    end
    endgenerate
    
    
    
    // LUT : 2019
    wire [63:0] lut_2019_table = 64'b0101010111011101010101011101010100000001100011010000000010000000;
    wire [5:0] lut_2019_select = {
                             in_data[351],
                             in_data[497],
                             in_data[399],
                             in_data[515],
                             in_data[522],
                             in_data[293]};
    
    wire lut_2019_out = lut_2019_table[lut_2019_select];
    
    generate
    if ( USE_REG ) begin : ff_2019
        reg   lut_2019_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2019_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2019_ff <= lut_2019_out;
            end
        end
        
        assign out_data[2019] = lut_2019_ff;
    end
    else begin : no_ff_2019
        assign out_data[2019] = lut_2019_out;
    end
    endgenerate
    
    
    
    // LUT : 2020
    wire [63:0] lut_2020_table = 64'b1101010001000000110000000000000011111111111111111111111011001100;
    wire [5:0] lut_2020_select = {
                             in_data[635],
                             in_data[545],
                             in_data[182],
                             in_data[193],
                             in_data[713],
                             in_data[533]};
    
    wire lut_2020_out = lut_2020_table[lut_2020_select];
    
    generate
    if ( USE_REG ) begin : ff_2020
        reg   lut_2020_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2020_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2020_ff <= lut_2020_out;
            end
        end
        
        assign out_data[2020] = lut_2020_ff;
    end
    else begin : no_ff_2020
        assign out_data[2020] = lut_2020_out;
    end
    endgenerate
    
    
    
    // LUT : 2021
    wire [63:0] lut_2021_table = 64'b1111111111111111000000001011111111111111111111110000000011001100;
    wire [5:0] lut_2021_select = {
                             in_data[133],
                             in_data[102],
                             in_data[312],
                             in_data[532],
                             in_data[649],
                             in_data[4]};
    
    wire lut_2021_out = lut_2021_table[lut_2021_select];
    
    generate
    if ( USE_REG ) begin : ff_2021
        reg   lut_2021_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2021_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2021_ff <= lut_2021_out;
            end
        end
        
        assign out_data[2021] = lut_2021_ff;
    end
    else begin : no_ff_2021
        assign out_data[2021] = lut_2021_out;
    end
    endgenerate
    
    
    
    // LUT : 2022
    wire [63:0] lut_2022_table = 64'b0000000010001100000011001000111100000000100010000000110011001111;
    wire [5:0] lut_2022_select = {
                             in_data[756],
                             in_data[680],
                             in_data[333],
                             in_data[682],
                             in_data[218],
                             in_data[502]};
    
    wire lut_2022_out = lut_2022_table[lut_2022_select];
    
    generate
    if ( USE_REG ) begin : ff_2022
        reg   lut_2022_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2022_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2022_ff <= lut_2022_out;
            end
        end
        
        assign out_data[2022] = lut_2022_ff;
    end
    else begin : no_ff_2022
        assign out_data[2022] = lut_2022_out;
    end
    endgenerate
    
    
    
    // LUT : 2023
    wire [63:0] lut_2023_table = 64'b0000000011000000000000001101000000000000010111110000000001011111;
    wire [5:0] lut_2023_select = {
                             in_data[463],
                             in_data[738],
                             in_data[329],
                             in_data[594],
                             in_data[548],
                             in_data[481]};
    
    wire lut_2023_out = lut_2023_table[lut_2023_select];
    
    generate
    if ( USE_REG ) begin : ff_2023
        reg   lut_2023_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2023_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2023_ff <= lut_2023_out;
            end
        end
        
        assign out_data[2023] = lut_2023_ff;
    end
    else begin : no_ff_2023
        assign out_data[2023] = lut_2023_out;
    end
    endgenerate
    
    
    
    // LUT : 2024
    wire [63:0] lut_2024_table = 64'b0000010000000011010101110111011100000000000000000000000000000011;
    wire [5:0] lut_2024_select = {
                             in_data[563],
                             in_data[302],
                             in_data[582],
                             in_data[650],
                             in_data[267],
                             in_data[688]};
    
    wire lut_2024_out = lut_2024_table[lut_2024_select];
    
    generate
    if ( USE_REG ) begin : ff_2024
        reg   lut_2024_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2024_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2024_ff <= lut_2024_out;
            end
        end
        
        assign out_data[2024] = lut_2024_ff;
    end
    else begin : no_ff_2024
        assign out_data[2024] = lut_2024_out;
    end
    endgenerate
    
    
    
    // LUT : 2025
    wire [63:0] lut_2025_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_2025_select = {
                             in_data[777],
                             in_data[550],
                             in_data[636],
                             in_data[163],
                             in_data[617],
                             in_data[698]};
    
    wire lut_2025_out = lut_2025_table[lut_2025_select];
    
    generate
    if ( USE_REG ) begin : ff_2025
        reg   lut_2025_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2025_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2025_ff <= lut_2025_out;
            end
        end
        
        assign out_data[2025] = lut_2025_ff;
    end
    else begin : no_ff_2025
        assign out_data[2025] = lut_2025_out;
    end
    endgenerate
    
    
    
    // LUT : 2026
    wire [63:0] lut_2026_table = 64'b0101010101010101000000000000000001010101010101010000000000000000;
    wire [5:0] lut_2026_select = {
                             in_data[755],
                             in_data[295],
                             in_data[140],
                             in_data[480],
                             in_data[143],
                             in_data[499]};
    
    wire lut_2026_out = lut_2026_table[lut_2026_select];
    
    generate
    if ( USE_REG ) begin : ff_2026
        reg   lut_2026_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2026_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2026_ff <= lut_2026_out;
            end
        end
        
        assign out_data[2026] = lut_2026_ff;
    end
    else begin : no_ff_2026
        assign out_data[2026] = lut_2026_out;
    end
    endgenerate
    
    
    
    // LUT : 2027
    wire [63:0] lut_2027_table = 64'b1001100110011011000100010001000100001001100110110000000100110011;
    wire [5:0] lut_2027_select = {
                             in_data[655],
                             in_data[130],
                             in_data[93],
                             in_data[417],
                             in_data[378],
                             in_data[461]};
    
    wire lut_2027_out = lut_2027_table[lut_2027_select];
    
    generate
    if ( USE_REG ) begin : ff_2027
        reg   lut_2027_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2027_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2027_ff <= lut_2027_out;
            end
        end
        
        assign out_data[2027] = lut_2027_ff;
    end
    else begin : no_ff_2027
        assign out_data[2027] = lut_2027_out;
    end
    endgenerate
    
    
    
    // LUT : 2028
    wire [63:0] lut_2028_table = 64'b1111111101111111111111110000000011111111000000001111111100000000;
    wire [5:0] lut_2028_select = {
                             in_data[641],
                             in_data[674],
                             in_data[210],
                             in_data[15],
                             in_data[394],
                             in_data[589]};
    
    wire lut_2028_out = lut_2028_table[lut_2028_select];
    
    generate
    if ( USE_REG ) begin : ff_2028
        reg   lut_2028_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2028_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2028_ff <= lut_2028_out;
            end
        end
        
        assign out_data[2028] = lut_2028_ff;
    end
    else begin : no_ff_2028
        assign out_data[2028] = lut_2028_out;
    end
    endgenerate
    
    
    
    // LUT : 2029
    wire [63:0] lut_2029_table = 64'b1111111111111111111111111111111101001111000011110100111100001111;
    wire [5:0] lut_2029_select = {
                             in_data[607],
                             in_data[58],
                             in_data[392],
                             in_data[268],
                             in_data[358],
                             in_data[622]};
    
    wire lut_2029_out = lut_2029_table[lut_2029_select];
    
    generate
    if ( USE_REG ) begin : ff_2029
        reg   lut_2029_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2029_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2029_ff <= lut_2029_out;
            end
        end
        
        assign out_data[2029] = lut_2029_ff;
    end
    else begin : no_ff_2029
        assign out_data[2029] = lut_2029_out;
    end
    endgenerate
    
    
    
    // LUT : 2030
    wire [63:0] lut_2030_table = 64'b0000000100000101111111111111111100000101000001010000010100000111;
    wire [5:0] lut_2030_select = {
                             in_data[386],
                             in_data[176],
                             in_data[31],
                             in_data[376],
                             in_data[87],
                             in_data[696]};
    
    wire lut_2030_out = lut_2030_table[lut_2030_select];
    
    generate
    if ( USE_REG ) begin : ff_2030
        reg   lut_2030_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2030_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2030_ff <= lut_2030_out;
            end
        end
        
        assign out_data[2030] = lut_2030_ff;
    end
    else begin : no_ff_2030
        assign out_data[2030] = lut_2030_out;
    end
    endgenerate
    
    
    
    // LUT : 2031
    wire [63:0] lut_2031_table = 64'b1100000011000000111001111100110111000000110000001100010111001111;
    wire [5:0] lut_2031_select = {
                             in_data[448],
                             in_data[297],
                             in_data[236],
                             in_data[346],
                             in_data[436],
                             in_data[728]};
    
    wire lut_2031_out = lut_2031_table[lut_2031_select];
    
    generate
    if ( USE_REG ) begin : ff_2031
        reg   lut_2031_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2031_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2031_ff <= lut_2031_out;
            end
        end
        
        assign out_data[2031] = lut_2031_ff;
    end
    else begin : no_ff_2031
        assign out_data[2031] = lut_2031_out;
    end
    endgenerate
    
    
    
    // LUT : 2032
    wire [63:0] lut_2032_table = 64'b1111111111111111000001000100010111011111110111010100000001000100;
    wire [5:0] lut_2032_select = {
                             in_data[776],
                             in_data[403],
                             in_data[752],
                             in_data[77],
                             in_data[677],
                             in_data[177]};
    
    wire lut_2032_out = lut_2032_table[lut_2032_select];
    
    generate
    if ( USE_REG ) begin : ff_2032
        reg   lut_2032_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2032_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2032_ff <= lut_2032_out;
            end
        end
        
        assign out_data[2032] = lut_2032_ff;
    end
    else begin : no_ff_2032
        assign out_data[2032] = lut_2032_out;
    end
    endgenerate
    
    
    
    // LUT : 2033
    wire [63:0] lut_2033_table = 64'b0000000000000000000000000010000010100000101000001010011110110101;
    wire [5:0] lut_2033_select = {
                             in_data[715],
                             in_data[466],
                             in_data[279],
                             in_data[317],
                             in_data[253],
                             in_data[653]};
    
    wire lut_2033_out = lut_2033_table[lut_2033_select];
    
    generate
    if ( USE_REG ) begin : ff_2033
        reg   lut_2033_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2033_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2033_ff <= lut_2033_out;
            end
        end
        
        assign out_data[2033] = lut_2033_ff;
    end
    else begin : no_ff_2033
        assign out_data[2033] = lut_2033_out;
    end
    endgenerate
    
    
    
    // LUT : 2034
    wire [63:0] lut_2034_table = 64'b1010101111111111101010101111111100000000001000100000000000000000;
    wire [5:0] lut_2034_select = {
                             in_data[600],
                             in_data[254],
                             in_data[353],
                             in_data[3],
                             in_data[531],
                             in_data[181]};
    
    wire lut_2034_out = lut_2034_table[lut_2034_select];
    
    generate
    if ( USE_REG ) begin : ff_2034
        reg   lut_2034_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2034_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2034_ff <= lut_2034_out;
            end
        end
        
        assign out_data[2034] = lut_2034_ff;
    end
    else begin : no_ff_2034
        assign out_data[2034] = lut_2034_out;
    end
    endgenerate
    
    
    
    // LUT : 2035
    wire [63:0] lut_2035_table = 64'b1000000011000100111111001100110010000000110001001111110011001100;
    wire [5:0] lut_2035_select = {
                             in_data[20],
                             in_data[284],
                             in_data[349],
                             in_data[191],
                             in_data[402],
                             in_data[624]};
    
    wire lut_2035_out = lut_2035_table[lut_2035_select];
    
    generate
    if ( USE_REG ) begin : ff_2035
        reg   lut_2035_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2035_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2035_ff <= lut_2035_out;
            end
        end
        
        assign out_data[2035] = lut_2035_ff;
    end
    else begin : no_ff_2035
        assign out_data[2035] = lut_2035_out;
    end
    endgenerate
    
    
    
    // LUT : 2036
    wire [63:0] lut_2036_table = 64'b1100000011000000111100001111000000000000000000001111000011110000;
    wire [5:0] lut_2036_select = {
                             in_data[774],
                             in_data[67],
                             in_data[561],
                             in_data[381],
                             in_data[382],
                             in_data[79]};
    
    wire lut_2036_out = lut_2036_table[lut_2036_select];
    
    generate
    if ( USE_REG ) begin : ff_2036
        reg   lut_2036_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2036_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2036_ff <= lut_2036_out;
            end
        end
        
        assign out_data[2036] = lut_2036_ff;
    end
    else begin : no_ff_2036
        assign out_data[2036] = lut_2036_out;
    end
    endgenerate
    
    
    
    // LUT : 2037
    wire [63:0] lut_2037_table = 64'b0101010101010101000000000000000001111111010101010101010101010000;
    wire [5:0] lut_2037_select = {
                             in_data[121],
                             in_data[256],
                             in_data[222],
                             in_data[471],
                             in_data[673],
                             in_data[719]};
    
    wire lut_2037_out = lut_2037_table[lut_2037_select];
    
    generate
    if ( USE_REG ) begin : ff_2037
        reg   lut_2037_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2037_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2037_ff <= lut_2037_out;
            end
        end
        
        assign out_data[2037] = lut_2037_ff;
    end
    else begin : no_ff_2037
        assign out_data[2037] = lut_2037_out;
    end
    endgenerate
    
    
    
    // LUT : 2038
    wire [63:0] lut_2038_table = 64'b1111111101010101000000000000000000010001010101010101010101010101;
    wire [5:0] lut_2038_select = {
                             in_data[187],
                             in_data[626],
                             in_data[741],
                             in_data[366],
                             in_data[106],
                             in_data[327]};
    
    wire lut_2038_out = lut_2038_table[lut_2038_select];
    
    generate
    if ( USE_REG ) begin : ff_2038
        reg   lut_2038_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2038_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2038_ff <= lut_2038_out;
            end
        end
        
        assign out_data[2038] = lut_2038_ff;
    end
    else begin : no_ff_2038
        assign out_data[2038] = lut_2038_out;
    end
    endgenerate
    
    
    
    // LUT : 2039
    wire [63:0] lut_2039_table = 64'b0100111111111111000000001111111100000000111111110000000000001111;
    wire [5:0] lut_2039_select = {
                             in_data[564],
                             in_data[200],
                             in_data[441],
                             in_data[446],
                             in_data[49],
                             in_data[419]};
    
    wire lut_2039_out = lut_2039_table[lut_2039_select];
    
    generate
    if ( USE_REG ) begin : ff_2039
        reg   lut_2039_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2039_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2039_ff <= lut_2039_out;
            end
        end
        
        assign out_data[2039] = lut_2039_ff;
    end
    else begin : no_ff_2039
        assign out_data[2039] = lut_2039_out;
    end
    endgenerate
    
    
    
    // LUT : 2040
    wire [63:0] lut_2040_table = 64'b0101010101010101010101010101010101010000010101010101000001010101;
    wire [5:0] lut_2040_select = {
                             in_data[492],
                             in_data[142],
                             in_data[258],
                             in_data[584],
                             in_data[420],
                             in_data[205]};
    
    wire lut_2040_out = lut_2040_table[lut_2040_select];
    
    generate
    if ( USE_REG ) begin : ff_2040
        reg   lut_2040_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2040_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2040_ff <= lut_2040_out;
            end
        end
        
        assign out_data[2040] = lut_2040_ff;
    end
    else begin : no_ff_2040
        assign out_data[2040] = lut_2040_out;
    end
    endgenerate
    
    
    
    // LUT : 2041
    wire [63:0] lut_2041_table = 64'b0000000010110011000000001111111100000000001100010000000011111111;
    wire [5:0] lut_2041_select = {
                             in_data[541],
                             in_data[483],
                             in_data[184],
                             in_data[169],
                             in_data[424],
                             in_data[726]};
    
    wire lut_2041_out = lut_2041_table[lut_2041_select];
    
    generate
    if ( USE_REG ) begin : ff_2041
        reg   lut_2041_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2041_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2041_ff <= lut_2041_out;
            end
        end
        
        assign out_data[2041] = lut_2041_ff;
    end
    else begin : no_ff_2041
        assign out_data[2041] = lut_2041_out;
    end
    endgenerate
    
    
    
    // LUT : 2042
    wire [63:0] lut_2042_table = 64'b1111111111111111000000001111111111111111111111110000000011111111;
    wire [5:0] lut_2042_select = {
                             in_data[697],
                             in_data[315],
                             in_data[185],
                             in_data[609],
                             in_data[36],
                             in_data[306]};
    
    wire lut_2042_out = lut_2042_table[lut_2042_select];
    
    generate
    if ( USE_REG ) begin : ff_2042
        reg   lut_2042_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2042_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2042_ff <= lut_2042_out;
            end
        end
        
        assign out_data[2042] = lut_2042_ff;
    end
    else begin : no_ff_2042
        assign out_data[2042] = lut_2042_out;
    end
    endgenerate
    
    
    
    // LUT : 2043
    wire [63:0] lut_2043_table = 64'b0101010101010101110111011101110101010101010101011101111111011101;
    wire [5:0] lut_2043_select = {
                             in_data[282],
                             in_data[457],
                             in_data[505],
                             in_data[88],
                             in_data[740],
                             in_data[577]};
    
    wire lut_2043_out = lut_2043_table[lut_2043_select];
    
    generate
    if ( USE_REG ) begin : ff_2043
        reg   lut_2043_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2043_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2043_ff <= lut_2043_out;
            end
        end
        
        assign out_data[2043] = lut_2043_ff;
    end
    else begin : no_ff_2043
        assign out_data[2043] = lut_2043_out;
    end
    endgenerate
    
    
    
    // LUT : 2044
    wire [63:0] lut_2044_table = 64'b1111111111111111111111111111111100001110000000000000111100001000;
    wire [5:0] lut_2044_select = {
                             in_data[491],
                             in_data[616],
                             in_data[519],
                             in_data[161],
                             in_data[575],
                             in_data[771]};
    
    wire lut_2044_out = lut_2044_table[lut_2044_select];
    
    generate
    if ( USE_REG ) begin : ff_2044
        reg   lut_2044_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2044_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2044_ff <= lut_2044_out;
            end
        end
        
        assign out_data[2044] = lut_2044_ff;
    end
    else begin : no_ff_2044
        assign out_data[2044] = lut_2044_out;
    end
    endgenerate
    
    
    
    // LUT : 2045
    wire [63:0] lut_2045_table = 64'b0000000000000000000000000000000000001010001100110000101000110011;
    wire [5:0] lut_2045_select = {
                             in_data[179],
                             in_data[197],
                             in_data[625],
                             in_data[334],
                             in_data[569],
                             in_data[25]};
    
    wire lut_2045_out = lut_2045_table[lut_2045_select];
    
    generate
    if ( USE_REG ) begin : ff_2045
        reg   lut_2045_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2045_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2045_ff <= lut_2045_out;
            end
        end
        
        assign out_data[2045] = lut_2045_ff;
    end
    else begin : no_ff_2045
        assign out_data[2045] = lut_2045_out;
    end
    endgenerate
    
    
    
    // LUT : 2046
    wire [63:0] lut_2046_table = 64'b0011001111111111001100111111111100110011111111110011001111101110;
    wire [5:0] lut_2046_select = {
                             in_data[782],
                             in_data[773],
                             in_data[454],
                             in_data[780],
                             in_data[345],
                             in_data[647]};
    
    wire lut_2046_out = lut_2046_table[lut_2046_select];
    
    generate
    if ( USE_REG ) begin : ff_2046
        reg   lut_2046_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2046_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2046_ff <= lut_2046_out;
            end
        end
        
        assign out_data[2046] = lut_2046_ff;
    end
    else begin : no_ff_2046
        assign out_data[2046] = lut_2046_out;
    end
    endgenerate
    
    
    
    // LUT : 2047
    wire [63:0] lut_2047_table = 64'b0000110000001100000011000000110010001111000011111110111100001111;
    wire [5:0] lut_2047_select = {
                             in_data[265],
                             in_data[587],
                             in_data[432],
                             in_data[209],
                             in_data[226],
                             in_data[590]};
    
    wire lut_2047_out = lut_2047_table[lut_2047_select];
    
    generate
    if ( USE_REG ) begin : ff_2047
        reg   lut_2047_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2047_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2047_ff <= lut_2047_out;
            end
        end
        
        assign out_data[2047] = lut_2047_ff;
    end
    else begin : no_ff_2047
        assign out_data[2047] = lut_2047_out;
    end
    endgenerate
    
    
    
    // LUT : 2048
    wire [63:0] lut_2048_table = 64'b1100111100001111110011110000111101001111000011110100111100001111;
    wire [5:0] lut_2048_select = {
                             in_data[654],
                             in_data[754],
                             in_data[231],
                             in_data[549],
                             in_data[521],
                             in_data[501]};
    
    wire lut_2048_out = lut_2048_table[lut_2048_select];
    
    generate
    if ( USE_REG ) begin : ff_2048
        reg   lut_2048_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2048_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2048_ff <= lut_2048_out;
            end
        end
        
        assign out_data[2048] = lut_2048_ff;
    end
    else begin : no_ff_2048
        assign out_data[2048] = lut_2048_out;
    end
    endgenerate
    
    
    
    // LUT : 2049
    wire [63:0] lut_2049_table = 64'b0000111100011111000000000000000000111111001111110000110000001100;
    wire [5:0] lut_2049_select = {
                             in_data[583],
                             in_data[320],
                             in_data[671],
                             in_data[634],
                             in_data[566],
                             in_data[35]};
    
    wire lut_2049_out = lut_2049_table[lut_2049_select];
    
    generate
    if ( USE_REG ) begin : ff_2049
        reg   lut_2049_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2049_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2049_ff <= lut_2049_out;
            end
        end
        
        assign out_data[2049] = lut_2049_ff;
    end
    else begin : no_ff_2049
        assign out_data[2049] = lut_2049_out;
    end
    endgenerate
    
    
    
    // LUT : 2050
    wire [63:0] lut_2050_table = 64'b0000000011001111000000001100111100000000110011110000000011001111;
    wire [5:0] lut_2050_select = {
                             in_data[52],
                             in_data[144],
                             in_data[573],
                             in_data[397],
                             in_data[708],
                             in_data[645]};
    
    wire lut_2050_out = lut_2050_table[lut_2050_select];
    
    generate
    if ( USE_REG ) begin : ff_2050
        reg   lut_2050_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2050_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2050_ff <= lut_2050_out;
            end
        end
        
        assign out_data[2050] = lut_2050_ff;
    end
    else begin : no_ff_2050
        assign out_data[2050] = lut_2050_out;
    end
    endgenerate
    
    
    
    // LUT : 2051
    wire [63:0] lut_2051_table = 64'b1111111111011111111111111101111011111111110111111111111000000000;
    wire [5:0] lut_2051_select = {
                             in_data[736],
                             in_data[459],
                             in_data[357],
                             in_data[275],
                             in_data[228],
                             in_data[547]};
    
    wire lut_2051_out = lut_2051_table[lut_2051_select];
    
    generate
    if ( USE_REG ) begin : ff_2051
        reg   lut_2051_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2051_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2051_ff <= lut_2051_out;
            end
        end
        
        assign out_data[2051] = lut_2051_ff;
    end
    else begin : no_ff_2051
        assign out_data[2051] = lut_2051_out;
    end
    endgenerate
    
    
    
    // LUT : 2052
    wire [63:0] lut_2052_table = 64'b1010101100000010101010110000001010101011000000100010101100000010;
    wire [5:0] lut_2052_select = {
                             in_data[37],
                             in_data[165],
                             in_data[552],
                             in_data[155],
                             in_data[415],
                             in_data[484]};
    
    wire lut_2052_out = lut_2052_table[lut_2052_select];
    
    generate
    if ( USE_REG ) begin : ff_2052
        reg   lut_2052_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2052_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2052_ff <= lut_2052_out;
            end
        end
        
        assign out_data[2052] = lut_2052_ff;
    end
    else begin : no_ff_2052
        assign out_data[2052] = lut_2052_out;
    end
    endgenerate
    
    
    
    // LUT : 2053
    wire [63:0] lut_2053_table = 64'b1110111011101110111011101110111011111111111111111110111011111111;
    wire [5:0] lut_2053_select = {
                             in_data[186],
                             in_data[455],
                             in_data[478],
                             in_data[81],
                             in_data[206],
                             in_data[303]};
    
    wire lut_2053_out = lut_2053_table[lut_2053_select];
    
    generate
    if ( USE_REG ) begin : ff_2053
        reg   lut_2053_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2053_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2053_ff <= lut_2053_out;
            end
        end
        
        assign out_data[2053] = lut_2053_ff;
    end
    else begin : no_ff_2053
        assign out_data[2053] = lut_2053_out;
    end
    endgenerate
    
    
    
    // LUT : 2054
    wire [63:0] lut_2054_table = 64'b0100010101010101000000000000000001010101010111110000000000000101;
    wire [5:0] lut_2054_select = {
                             in_data[724],
                             in_data[194],
                             in_data[118],
                             in_data[389],
                             in_data[60],
                             in_data[444]};
    
    wire lut_2054_out = lut_2054_table[lut_2054_select];
    
    generate
    if ( USE_REG ) begin : ff_2054
        reg   lut_2054_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2054_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2054_ff <= lut_2054_out;
            end
        end
        
        assign out_data[2054] = lut_2054_ff;
    end
    else begin : no_ff_2054
        assign out_data[2054] = lut_2054_out;
    end
    endgenerate
    
    
    
    // LUT : 2055
    wire [63:0] lut_2055_table = 64'b1011101110111011101010111011101110111011101110111011101110111011;
    wire [5:0] lut_2055_select = {
                             in_data[758],
                             in_data[721],
                             in_data[685],
                             in_data[30],
                             in_data[604],
                             in_data[369]};
    
    wire lut_2055_out = lut_2055_table[lut_2055_select];
    
    generate
    if ( USE_REG ) begin : ff_2055
        reg   lut_2055_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2055_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2055_ff <= lut_2055_out;
            end
        end
        
        assign out_data[2055] = lut_2055_ff;
    end
    else begin : no_ff_2055
        assign out_data[2055] = lut_2055_out;
    end
    endgenerate
    
    
    
    // LUT : 2056
    wire [63:0] lut_2056_table = 64'b1110111111001100111111111111111111001101000000001100110001000100;
    wire [5:0] lut_2056_select = {
                             in_data[404],
                             in_data[469],
                             in_data[570],
                             in_data[11],
                             in_data[665],
                             in_data[712]};
    
    wire lut_2056_out = lut_2056_table[lut_2056_select];
    
    generate
    if ( USE_REG ) begin : ff_2056
        reg   lut_2056_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2056_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2056_ff <= lut_2056_out;
            end
        end
        
        assign out_data[2056] = lut_2056_ff;
    end
    else begin : no_ff_2056
        assign out_data[2056] = lut_2056_out;
    end
    endgenerate
    
    
    
    // LUT : 2057
    wire [63:0] lut_2057_table = 64'b0000111111111111000011111110111111001111111111111100110011001100;
    wire [5:0] lut_2057_select = {
                             in_data[512],
                             in_data[578],
                             in_data[375],
                             in_data[242],
                             in_data[538],
                             in_data[195]};
    
    wire lut_2057_out = lut_2057_table[lut_2057_select];
    
    generate
    if ( USE_REG ) begin : ff_2057
        reg   lut_2057_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2057_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2057_ff <= lut_2057_out;
            end
        end
        
        assign out_data[2057] = lut_2057_ff;
    end
    else begin : no_ff_2057
        assign out_data[2057] = lut_2057_out;
    end
    endgenerate
    
    
    
    // LUT : 2058
    wire [63:0] lut_2058_table = 64'b1100110011001100110011001100110011001101110011000000110001001100;
    wire [5:0] lut_2058_select = {
                             in_data[154],
                             in_data[380],
                             in_data[304],
                             in_data[681],
                             in_data[264],
                             in_data[722]};
    
    wire lut_2058_out = lut_2058_table[lut_2058_select];
    
    generate
    if ( USE_REG ) begin : ff_2058
        reg   lut_2058_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2058_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2058_ff <= lut_2058_out;
            end
        end
        
        assign out_data[2058] = lut_2058_ff;
    end
    else begin : no_ff_2058
        assign out_data[2058] = lut_2058_out;
    end
    endgenerate
    
    
    
    // LUT : 2059
    wire [63:0] lut_2059_table = 64'b1111111111111111110011111100111111001111110011111000111110001100;
    wire [5:0] lut_2059_select = {
                             in_data[396],
                             in_data[368],
                             in_data[14],
                             in_data[180],
                             in_data[438],
                             in_data[63]};
    
    wire lut_2059_out = lut_2059_table[lut_2059_select];
    
    generate
    if ( USE_REG ) begin : ff_2059
        reg   lut_2059_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2059_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2059_ff <= lut_2059_out;
            end
        end
        
        assign out_data[2059] = lut_2059_ff;
    end
    else begin : no_ff_2059
        assign out_data[2059] = lut_2059_out;
    end
    endgenerate
    
    
    
    // LUT : 2060
    wire [63:0] lut_2060_table = 64'b1100010011110000111010111111111111000000110000001110100011111111;
    wire [5:0] lut_2060_select = {
                             in_data[227],
                             in_data[660],
                             in_data[692],
                             in_data[716],
                             in_data[453],
                             in_data[245]};
    
    wire lut_2060_out = lut_2060_table[lut_2060_select];
    
    generate
    if ( USE_REG ) begin : ff_2060
        reg   lut_2060_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2060_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2060_ff <= lut_2060_out;
            end
        end
        
        assign out_data[2060] = lut_2060_ff;
    end
    else begin : no_ff_2060
        assign out_data[2060] = lut_2060_out;
    end
    endgenerate
    
    
    
    // LUT : 2061
    wire [63:0] lut_2061_table = 64'b1111000000010000111110111101000011110000010100001111111111110000;
    wire [5:0] lut_2061_select = {
                             in_data[86],
                             in_data[526],
                             in_data[373],
                             in_data[629],
                             in_data[439],
                             in_data[460]};
    
    wire lut_2061_out = lut_2061_table[lut_2061_select];
    
    generate
    if ( USE_REG ) begin : ff_2061
        reg   lut_2061_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2061_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2061_ff <= lut_2061_out;
            end
        end
        
        assign out_data[2061] = lut_2061_ff;
    end
    else begin : no_ff_2061
        assign out_data[2061] = lut_2061_out;
    end
    endgenerate
    
    
    
    // LUT : 2062
    wire [63:0] lut_2062_table = 64'b1111000011110000111100111111001011110000111100001111001011110010;
    wire [5:0] lut_2062_select = {
                             in_data[672],
                             in_data[157],
                             in_data[69],
                             in_data[576],
                             in_data[518],
                             in_data[395]};
    
    wire lut_2062_out = lut_2062_table[lut_2062_select];
    
    generate
    if ( USE_REG ) begin : ff_2062
        reg   lut_2062_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2062_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2062_ff <= lut_2062_out;
            end
        end
        
        assign out_data[2062] = lut_2062_ff;
    end
    else begin : no_ff_2062
        assign out_data[2062] = lut_2062_out;
    end
    endgenerate
    
    
    
    // LUT : 2063
    wire [63:0] lut_2063_table = 64'b0001000011111111001000001111111100000000111100100000000011110011;
    wire [5:0] lut_2063_select = {
                             in_data[183],
                             in_data[477],
                             in_data[458],
                             in_data[678],
                             in_data[135],
                             in_data[19]};
    
    wire lut_2063_out = lut_2063_table[lut_2063_select];
    
    generate
    if ( USE_REG ) begin : ff_2063
        reg   lut_2063_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2063_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2063_ff <= lut_2063_out;
            end
        end
        
        assign out_data[2063] = lut_2063_ff;
    end
    else begin : no_ff_2063
        assign out_data[2063] = lut_2063_out;
    end
    endgenerate
    
    
    
    // LUT : 2064
    wire [63:0] lut_2064_table = 64'b0000000000000000000000000000000000000000010101010000000001010001;
    wire [5:0] lut_2064_select = {
                             in_data[534],
                             in_data[670],
                             in_data[612],
                             in_data[762],
                             in_data[115],
                             in_data[219]};
    
    wire lut_2064_out = lut_2064_table[lut_2064_select];
    
    generate
    if ( USE_REG ) begin : ff_2064
        reg   lut_2064_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2064_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2064_ff <= lut_2064_out;
            end
        end
        
        assign out_data[2064] = lut_2064_ff;
    end
    else begin : no_ff_2064
        assign out_data[2064] = lut_2064_out;
    end
    endgenerate
    
    
    
    // LUT : 2065
    wire [63:0] lut_2065_table = 64'b1111000011110000111100001111000011110011111100111111001111110011;
    wire [5:0] lut_2065_select = {
                             in_data[126],
                             in_data[278],
                             in_data[648],
                             in_data[658],
                             in_data[524],
                             in_data[2]};
    
    wire lut_2065_out = lut_2065_table[lut_2065_select];
    
    generate
    if ( USE_REG ) begin : ff_2065
        reg   lut_2065_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2065_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2065_ff <= lut_2065_out;
            end
        end
        
        assign out_data[2065] = lut_2065_ff;
    end
    else begin : no_ff_2065
        assign out_data[2065] = lut_2065_out;
    end
    endgenerate
    
    
    
    // LUT : 2066
    wire [63:0] lut_2066_table = 64'b1111111100000000111111110000000011111111111100001111111110100000;
    wire [5:0] lut_2066_select = {
                             in_data[137],
                             in_data[729],
                             in_data[398],
                             in_data[435],
                             in_data[251],
                             in_data[336]};
    
    wire lut_2066_out = lut_2066_table[lut_2066_select];
    
    generate
    if ( USE_REG ) begin : ff_2066
        reg   lut_2066_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2066_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2066_ff <= lut_2066_out;
            end
        end
        
        assign out_data[2066] = lut_2066_ff;
    end
    else begin : no_ff_2066
        assign out_data[2066] = lut_2066_out;
    end
    endgenerate
    
    
    
    // LUT : 2067
    wire [63:0] lut_2067_table = 64'b1111111111111111001100110011001011111111111111110011001100000000;
    wire [5:0] lut_2067_select = {
                             in_data[472],
                             in_data[400],
                             in_data[414],
                             in_data[586],
                             in_data[652],
                             in_data[750]};
    
    wire lut_2067_out = lut_2067_table[lut_2067_select];
    
    generate
    if ( USE_REG ) begin : ff_2067
        reg   lut_2067_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2067_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2067_ff <= lut_2067_out;
            end
        end
        
        assign out_data[2067] = lut_2067_ff;
    end
    else begin : no_ff_2067
        assign out_data[2067] = lut_2067_out;
    end
    endgenerate
    
    
    
    // LUT : 2068
    wire [63:0] lut_2068_table = 64'b1011111100101111101111110010101110111111000010110011111100001111;
    wire [5:0] lut_2068_select = {
                             in_data[73],
                             in_data[281],
                             in_data[510],
                             in_data[409],
                             in_data[428],
                             in_data[237]};
    
    wire lut_2068_out = lut_2068_table[lut_2068_select];
    
    generate
    if ( USE_REG ) begin : ff_2068
        reg   lut_2068_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2068_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2068_ff <= lut_2068_out;
            end
        end
        
        assign out_data[2068] = lut_2068_ff;
    end
    else begin : no_ff_2068
        assign out_data[2068] = lut_2068_out;
    end
    endgenerate
    
    
    
    // LUT : 2069
    wire [63:0] lut_2069_table = 64'b1111111111111111111111111111111111111111000010001111111100000000;
    wire [5:0] lut_2069_select = {
                             in_data[216],
                             in_data[170],
                             in_data[487],
                             in_data[319],
                             in_data[41],
                             in_data[252]};
    
    wire lut_2069_out = lut_2069_table[lut_2069_select];
    
    generate
    if ( USE_REG ) begin : ff_2069
        reg   lut_2069_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2069_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2069_ff <= lut_2069_out;
            end
        end
        
        assign out_data[2069] = lut_2069_ff;
    end
    else begin : no_ff_2069
        assign out_data[2069] = lut_2069_out;
    end
    endgenerate
    
    
    
    // LUT : 2070
    wire [63:0] lut_2070_table = 64'b1111010110100101111101011010010111110101000001000001010100000100;
    wire [5:0] lut_2070_select = {
                             in_data[711],
                             in_data[763],
                             in_data[599],
                             in_data[271],
                             in_data[43],
                             in_data[244]};
    
    wire lut_2070_out = lut_2070_table[lut_2070_select];
    
    generate
    if ( USE_REG ) begin : ff_2070
        reg   lut_2070_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2070_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2070_ff <= lut_2070_out;
            end
        end
        
        assign out_data[2070] = lut_2070_ff;
    end
    else begin : no_ff_2070
        assign out_data[2070] = lut_2070_out;
    end
    endgenerate
    
    
    
    // LUT : 2071
    wire [63:0] lut_2071_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_2071_select = {
                             in_data[116],
                             in_data[579],
                             in_data[298],
                             in_data[707],
                             in_data[110],
                             in_data[199]};
    
    wire lut_2071_out = lut_2071_table[lut_2071_select];
    
    generate
    if ( USE_REG ) begin : ff_2071
        reg   lut_2071_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2071_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2071_ff <= lut_2071_out;
            end
        end
        
        assign out_data[2071] = lut_2071_ff;
    end
    else begin : no_ff_2071
        assign out_data[2071] = lut_2071_out;
    end
    endgenerate
    
    
    
    // LUT : 2072
    wire [63:0] lut_2072_table = 64'b0000111100001111000010000000000011101111101011111111111111111111;
    wire [5:0] lut_2072_select = {
                             in_data[407],
                             in_data[493],
                             in_data[223],
                             in_data[508],
                             in_data[644],
                             in_data[694]};
    
    wire lut_2072_out = lut_2072_table[lut_2072_select];
    
    generate
    if ( USE_REG ) begin : ff_2072
        reg   lut_2072_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2072_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2072_ff <= lut_2072_out;
            end
        end
        
        assign out_data[2072] = lut_2072_ff;
    end
    else begin : no_ff_2072
        assign out_data[2072] = lut_2072_out;
    end
    endgenerate
    
    
    
    // LUT : 2073
    wire [63:0] lut_2073_table = 64'b0101010101010101010101010101010100000000000000000000000000000000;
    wire [5:0] lut_2073_select = {
                             in_data[430],
                             in_data[580],
                             in_data[775],
                             in_data[249],
                             in_data[702],
                             in_data[148]};
    
    wire lut_2073_out = lut_2073_table[lut_2073_select];
    
    generate
    if ( USE_REG ) begin : ff_2073
        reg   lut_2073_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2073_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2073_ff <= lut_2073_out;
            end
        end
        
        assign out_data[2073] = lut_2073_ff;
    end
    else begin : no_ff_2073
        assign out_data[2073] = lut_2073_out;
    end
    endgenerate
    
    
    
    // LUT : 2074
    wire [63:0] lut_2074_table = 64'b0000010100001101000001010000110100000101000011010000010100001101;
    wire [5:0] lut_2074_select = {
                             in_data[17],
                             in_data[114],
                             in_data[196],
                             in_data[44],
                             in_data[768],
                             in_data[356]};
    
    wire lut_2074_out = lut_2074_table[lut_2074_select];
    
    generate
    if ( USE_REG ) begin : ff_2074
        reg   lut_2074_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2074_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2074_ff <= lut_2074_out;
            end
        end
        
        assign out_data[2074] = lut_2074_ff;
    end
    else begin : no_ff_2074
        assign out_data[2074] = lut_2074_out;
    end
    endgenerate
    
    
    
    // LUT : 2075
    wire [63:0] lut_2075_table = 64'b0000000000000000111111111111111100000000000000001111111111111111;
    wire [5:0] lut_2075_select = {
                             in_data[26],
                             in_data[514],
                             in_data[760],
                             in_data[498],
                             in_data[296],
                             in_data[723]};
    
    wire lut_2075_out = lut_2075_table[lut_2075_select];
    
    generate
    if ( USE_REG ) begin : ff_2075
        reg   lut_2075_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2075_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2075_ff <= lut_2075_out;
            end
        end
        
        assign out_data[2075] = lut_2075_ff;
    end
    else begin : no_ff_2075
        assign out_data[2075] = lut_2075_out;
    end
    endgenerate
    
    
    
    // LUT : 2076
    wire [63:0] lut_2076_table = 64'b1011101010111111101010101010101010111011111111111010101010111111;
    wire [5:0] lut_2076_select = {
                             in_data[535],
                             in_data[684],
                             in_data[408],
                             in_data[744],
                             in_data[772],
                             in_data[662]};
    
    wire lut_2076_out = lut_2076_table[lut_2076_select];
    
    generate
    if ( USE_REG ) begin : ff_2076
        reg   lut_2076_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2076_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2076_ff <= lut_2076_out;
            end
        end
        
        assign out_data[2076] = lut_2076_ff;
    end
    else begin : no_ff_2076
        assign out_data[2076] = lut_2076_out;
    end
    endgenerate
    
    
    
    // LUT : 2077
    wire [63:0] lut_2077_table = 64'b0000000011111111000000001111111110100000111111110000000011111111;
    wire [5:0] lut_2077_select = {
                             in_data[468],
                             in_data[679],
                             in_data[238],
                             in_data[543],
                             in_data[56],
                             in_data[393]};
    
    wire lut_2077_out = lut_2077_table[lut_2077_select];
    
    generate
    if ( USE_REG ) begin : ff_2077
        reg   lut_2077_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2077_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2077_ff <= lut_2077_out;
            end
        end
        
        assign out_data[2077] = lut_2077_ff;
    end
    else begin : no_ff_2077
        assign out_data[2077] = lut_2077_out;
    end
    endgenerate
    
    
    
    // LUT : 2078
    wire [63:0] lut_2078_table = 64'b0011111100111111000000000000000000111111001111110000000000000000;
    wire [5:0] lut_2078_select = {
                             in_data[562],
                             in_data[627],
                             in_data[225],
                             in_data[212],
                             in_data[689],
                             in_data[618]};
    
    wire lut_2078_out = lut_2078_table[lut_2078_select];
    
    generate
    if ( USE_REG ) begin : ff_2078
        reg   lut_2078_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2078_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2078_ff <= lut_2078_out;
            end
        end
        
        assign out_data[2078] = lut_2078_ff;
    end
    else begin : no_ff_2078
        assign out_data[2078] = lut_2078_out;
    end
    endgenerate
    
    
    
    // LUT : 2079
    wire [63:0] lut_2079_table = 64'b1110111011001100110011101100110011111111111011101111111111101110;
    wire [5:0] lut_2079_select = {
                             in_data[305],
                             in_data[111],
                             in_data[717],
                             in_data[596],
                             in_data[202],
                             in_data[91]};
    
    wire lut_2079_out = lut_2079_table[lut_2079_select];
    
    generate
    if ( USE_REG ) begin : ff_2079
        reg   lut_2079_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2079_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2079_ff <= lut_2079_out;
            end
        end
        
        assign out_data[2079] = lut_2079_ff;
    end
    else begin : no_ff_2079
        assign out_data[2079] = lut_2079_out;
    end
    endgenerate
    
    
    
    // LUT : 2080
    wire [63:0] lut_2080_table = 64'b0000000010110011000000000011001000000010111100110000001010110011;
    wire [5:0] lut_2080_select = {
                             in_data[766],
                             in_data[754],
                             in_data[593],
                             in_data[412],
                             in_data[657],
                             in_data[98]};
    
    wire lut_2080_out = lut_2080_table[lut_2080_select];
    
    generate
    if ( USE_REG ) begin : ff_2080
        reg   lut_2080_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2080_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2080_ff <= lut_2080_out;
            end
        end
        
        assign out_data[2080] = lut_2080_ff;
    end
    else begin : no_ff_2080
        assign out_data[2080] = lut_2080_out;
    end
    endgenerate
    
    
    
    // LUT : 2081
    wire [63:0] lut_2081_table = 64'b0011001100111111001100111111111100110011001111110011001100111111;
    wire [5:0] lut_2081_select = {
                             in_data[506],
                             in_data[45],
                             in_data[372],
                             in_data[20],
                             in_data[410],
                             in_data[54]};
    
    wire lut_2081_out = lut_2081_table[lut_2081_select];
    
    generate
    if ( USE_REG ) begin : ff_2081
        reg   lut_2081_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2081_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2081_ff <= lut_2081_out;
            end
        end
        
        assign out_data[2081] = lut_2081_ff;
    end
    else begin : no_ff_2081
        assign out_data[2081] = lut_2081_out;
    end
    endgenerate
    
    
    
    // LUT : 2082
    wire [63:0] lut_2082_table = 64'b0000000000000000111011111100111000000000000000001111111111001110;
    wire [5:0] lut_2082_select = {
                             in_data[759],
                             in_data[303],
                             in_data[10],
                             in_data[775],
                             in_data[99],
                             in_data[41]};
    
    wire lut_2082_out = lut_2082_table[lut_2082_select];
    
    generate
    if ( USE_REG ) begin : ff_2082
        reg   lut_2082_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2082_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2082_ff <= lut_2082_out;
            end
        end
        
        assign out_data[2082] = lut_2082_ff;
    end
    else begin : no_ff_2082
        assign out_data[2082] = lut_2082_out;
    end
    endgenerate
    
    
    
    // LUT : 2083
    wire [63:0] lut_2083_table = 64'b1100110011001100111111111111111111001100110011001111111111111111;
    wire [5:0] lut_2083_select = {
                             in_data[612],
                             in_data[343],
                             in_data[138],
                             in_data[774],
                             in_data[536],
                             in_data[61]};
    
    wire lut_2083_out = lut_2083_table[lut_2083_select];
    
    generate
    if ( USE_REG ) begin : ff_2083
        reg   lut_2083_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2083_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2083_ff <= lut_2083_out;
            end
        end
        
        assign out_data[2083] = lut_2083_ff;
    end
    else begin : no_ff_2083
        assign out_data[2083] = lut_2083_out;
    end
    endgenerate
    
    
    
    // LUT : 2084
    wire [63:0] lut_2084_table = 64'b1111111110110010111111111011001011111111101100101111111110110010;
    wire [5:0] lut_2084_select = {
                             in_data[142],
                             in_data[670],
                             in_data[443],
                             in_data[737],
                             in_data[332],
                             in_data[257]};
    
    wire lut_2084_out = lut_2084_table[lut_2084_select];
    
    generate
    if ( USE_REG ) begin : ff_2084
        reg   lut_2084_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2084_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2084_ff <= lut_2084_out;
            end
        end
        
        assign out_data[2084] = lut_2084_ff;
    end
    else begin : no_ff_2084
        assign out_data[2084] = lut_2084_out;
    end
    endgenerate
    
    
    
    // LUT : 2085
    wire [63:0] lut_2085_table = 64'b1100110000000000110011001100110011001100110011001100110111011100;
    wire [5:0] lut_2085_select = {
                             in_data[316],
                             in_data[738],
                             in_data[156],
                             in_data[724],
                             in_data[326],
                             in_data[632]};
    
    wire lut_2085_out = lut_2085_table[lut_2085_select];
    
    generate
    if ( USE_REG ) begin : ff_2085
        reg   lut_2085_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2085_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2085_ff <= lut_2085_out;
            end
        end
        
        assign out_data[2085] = lut_2085_ff;
    end
    else begin : no_ff_2085
        assign out_data[2085] = lut_2085_out;
    end
    endgenerate
    
    
    
    // LUT : 2086
    wire [63:0] lut_2086_table = 64'b0000000000000000000000000000000011001100110011111100110011001111;
    wire [5:0] lut_2086_select = {
                             in_data[271],
                             in_data[140],
                             in_data[208],
                             in_data[607],
                             in_data[189],
                             in_data[673]};
    
    wire lut_2086_out = lut_2086_table[lut_2086_select];
    
    generate
    if ( USE_REG ) begin : ff_2086
        reg   lut_2086_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2086_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2086_ff <= lut_2086_out;
            end
        end
        
        assign out_data[2086] = lut_2086_ff;
    end
    else begin : no_ff_2086
        assign out_data[2086] = lut_2086_out;
    end
    endgenerate
    
    
    
    // LUT : 2087
    wire [63:0] lut_2087_table = 64'b1100100011001100110111001101110011000000110011001101110011011100;
    wire [5:0] lut_2087_select = {
                             in_data[717],
                             in_data[716],
                             in_data[720],
                             in_data[77],
                             in_data[371],
                             in_data[174]};
    
    wire lut_2087_out = lut_2087_table[lut_2087_select];
    
    generate
    if ( USE_REG ) begin : ff_2087
        reg   lut_2087_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2087_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2087_ff <= lut_2087_out;
            end
        end
        
        assign out_data[2087] = lut_2087_ff;
    end
    else begin : no_ff_2087
        assign out_data[2087] = lut_2087_out;
    end
    endgenerate
    
    
    
    // LUT : 2088
    wire [63:0] lut_2088_table = 64'b0000000000000000000000000000111000001000000011000000111000001100;
    wire [5:0] lut_2088_select = {
                             in_data[538],
                             in_data[479],
                             in_data[329],
                             in_data[556],
                             in_data[429],
                             in_data[772]};
    
    wire lut_2088_out = lut_2088_table[lut_2088_select];
    
    generate
    if ( USE_REG ) begin : ff_2088
        reg   lut_2088_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2088_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2088_ff <= lut_2088_out;
            end
        end
        
        assign out_data[2088] = lut_2088_ff;
    end
    else begin : no_ff_2088
        assign out_data[2088] = lut_2088_out;
    end
    endgenerate
    
    
    
    // LUT : 2089
    wire [63:0] lut_2089_table = 64'b0000000000001101000000000000110100000000000011110000000000001101;
    wire [5:0] lut_2089_select = {
                             in_data[113],
                             in_data[336],
                             in_data[76],
                             in_data[379],
                             in_data[734],
                             in_data[565]};
    
    wire lut_2089_out = lut_2089_table[lut_2089_select];
    
    generate
    if ( USE_REG ) begin : ff_2089
        reg   lut_2089_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2089_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2089_ff <= lut_2089_out;
            end
        end
        
        assign out_data[2089] = lut_2089_ff;
    end
    else begin : no_ff_2089
        assign out_data[2089] = lut_2089_out;
    end
    endgenerate
    
    
    
    // LUT : 2090
    wire [63:0] lut_2090_table = 64'b0101000001010000011100000111000001010100010101000101000001010000;
    wire [5:0] lut_2090_select = {
                             in_data[456],
                             in_data[596],
                             in_data[760],
                             in_data[237],
                             in_data[621],
                             in_data[512]};
    
    wire lut_2090_out = lut_2090_table[lut_2090_select];
    
    generate
    if ( USE_REG ) begin : ff_2090
        reg   lut_2090_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2090_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2090_ff <= lut_2090_out;
            end
        end
        
        assign out_data[2090] = lut_2090_ff;
    end
    else begin : no_ff_2090
        assign out_data[2090] = lut_2090_out;
    end
    endgenerate
    
    
    
    // LUT : 2091
    wire [63:0] lut_2091_table = 64'b1111111111111111111111001111110011111111111111111111110011111100;
    wire [5:0] lut_2091_select = {
                             in_data[503],
                             in_data[463],
                             in_data[82],
                             in_data[651],
                             in_data[460],
                             in_data[27]};
    
    wire lut_2091_out = lut_2091_table[lut_2091_select];
    
    generate
    if ( USE_REG ) begin : ff_2091
        reg   lut_2091_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2091_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2091_ff <= lut_2091_out;
            end
        end
        
        assign out_data[2091] = lut_2091_ff;
    end
    else begin : no_ff_2091
        assign out_data[2091] = lut_2091_out;
    end
    endgenerate
    
    
    
    // LUT : 2092
    wire [63:0] lut_2092_table = 64'b0001000100110011000000000000000000010001001100110000000000000000;
    wire [5:0] lut_2092_select = {
                             in_data[614],
                             in_data[294],
                             in_data[423],
                             in_data[730],
                             in_data[149],
                             in_data[171]};
    
    wire lut_2092_out = lut_2092_table[lut_2092_select];
    
    generate
    if ( USE_REG ) begin : ff_2092
        reg   lut_2092_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2092_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2092_ff <= lut_2092_out;
            end
        end
        
        assign out_data[2092] = lut_2092_ff;
    end
    else begin : no_ff_2092
        assign out_data[2092] = lut_2092_out;
    end
    endgenerate
    
    
    
    // LUT : 2093
    wire [63:0] lut_2093_table = 64'b0011001100110011001100110011001000110011001100110011001100110000;
    wire [5:0] lut_2093_select = {
                             in_data[64],
                             in_data[488],
                             in_data[388],
                             in_data[665],
                             in_data[592],
                             in_data[65]};
    
    wire lut_2093_out = lut_2093_table[lut_2093_select];
    
    generate
    if ( USE_REG ) begin : ff_2093
        reg   lut_2093_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2093_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2093_ff <= lut_2093_out;
            end
        end
        
        assign out_data[2093] = lut_2093_ff;
    end
    else begin : no_ff_2093
        assign out_data[2093] = lut_2093_out;
    end
    endgenerate
    
    
    
    // LUT : 2094
    wire [63:0] lut_2094_table = 64'b1111111111111111000000001111110011111101111111110000000011000000;
    wire [5:0] lut_2094_select = {
                             in_data[499],
                             in_data[295],
                             in_data[260],
                             in_data[546],
                             in_data[563],
                             in_data[193]};
    
    wire lut_2094_out = lut_2094_table[lut_2094_select];
    
    generate
    if ( USE_REG ) begin : ff_2094
        reg   lut_2094_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2094_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2094_ff <= lut_2094_out;
            end
        end
        
        assign out_data[2094] = lut_2094_ff;
    end
    else begin : no_ff_2094
        assign out_data[2094] = lut_2094_out;
    end
    endgenerate
    
    
    
    // LUT : 2095
    wire [63:0] lut_2095_table = 64'b0000000000000000000000000000000000000000001100110000000000110011;
    wire [5:0] lut_2095_select = {
                             in_data[267],
                             in_data[38],
                             in_data[321],
                             in_data[700],
                             in_data[191],
                             in_data[701]};
    
    wire lut_2095_out = lut_2095_table[lut_2095_select];
    
    generate
    if ( USE_REG ) begin : ff_2095
        reg   lut_2095_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2095_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2095_ff <= lut_2095_out;
            end
        end
        
        assign out_data[2095] = lut_2095_ff;
    end
    else begin : no_ff_2095
        assign out_data[2095] = lut_2095_out;
    end
    endgenerate
    
    
    
    // LUT : 2096
    wire [63:0] lut_2096_table = 64'b0000111100011111000010110000101100000111000001010000000000000000;
    wire [5:0] lut_2096_select = {
                             in_data[213],
                             in_data[510],
                             in_data[703],
                             in_data[441],
                             in_data[105],
                             in_data[302]};
    
    wire lut_2096_out = lut_2096_table[lut_2096_select];
    
    generate
    if ( USE_REG ) begin : ff_2096
        reg   lut_2096_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2096_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2096_ff <= lut_2096_out;
            end
        end
        
        assign out_data[2096] = lut_2096_ff;
    end
    else begin : no_ff_2096
        assign out_data[2096] = lut_2096_out;
    end
    endgenerate
    
    
    
    // LUT : 2097
    wire [63:0] lut_2097_table = 64'b0101000001010000010100000101000001010000010100000101000001010000;
    wire [5:0] lut_2097_select = {
                             in_data[420],
                             in_data[100],
                             in_data[196],
                             in_data[655],
                             in_data[29],
                             in_data[582]};
    
    wire lut_2097_out = lut_2097_table[lut_2097_select];
    
    generate
    if ( USE_REG ) begin : ff_2097
        reg   lut_2097_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2097_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2097_ff <= lut_2097_out;
            end
        end
        
        assign out_data[2097] = lut_2097_ff;
    end
    else begin : no_ff_2097
        assign out_data[2097] = lut_2097_out;
    end
    endgenerate
    
    
    
    // LUT : 2098
    wire [63:0] lut_2098_table = 64'b0000000000000000000000001111111100000000000000000000000011111111;
    wire [5:0] lut_2098_select = {
                             in_data[354],
                             in_data[468],
                             in_data[666],
                             in_data[714],
                             in_data[252],
                             in_data[782]};
    
    wire lut_2098_out = lut_2098_table[lut_2098_select];
    
    generate
    if ( USE_REG ) begin : ff_2098
        reg   lut_2098_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2098_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2098_ff <= lut_2098_out;
            end
        end
        
        assign out_data[2098] = lut_2098_ff;
    end
    else begin : no_ff_2098
        assign out_data[2098] = lut_2098_out;
    end
    endgenerate
    
    
    
    // LUT : 2099
    wire [63:0] lut_2099_table = 64'b1011111111111111000000000000000011111111101111110000000000000000;
    wire [5:0] lut_2099_select = {
                             in_data[606],
                             in_data[598],
                             in_data[139],
                             in_data[529],
                             in_data[301],
                             in_data[35]};
    
    wire lut_2099_out = lut_2099_table[lut_2099_select];
    
    generate
    if ( USE_REG ) begin : ff_2099
        reg   lut_2099_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2099_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2099_ff <= lut_2099_out;
            end
        end
        
        assign out_data[2099] = lut_2099_ff;
    end
    else begin : no_ff_2099
        assign out_data[2099] = lut_2099_out;
    end
    endgenerate
    
    
    
    // LUT : 2100
    wire [63:0] lut_2100_table = 64'b1100110011001100110011001100110011101111111111111110111111111111;
    wire [5:0] lut_2100_select = {
                             in_data[465],
                             in_data[16],
                             in_data[31],
                             in_data[781],
                             in_data[578],
                             in_data[531]};
    
    wire lut_2100_out = lut_2100_table[lut_2100_select];
    
    generate
    if ( USE_REG ) begin : ff_2100
        reg   lut_2100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2100_ff <= lut_2100_out;
            end
        end
        
        assign out_data[2100] = lut_2100_ff;
    end
    else begin : no_ff_2100
        assign out_data[2100] = lut_2100_out;
    end
    endgenerate
    
    
    
    // LUT : 2101
    wire [63:0] lut_2101_table = 64'b1011111100000000000011110000000000000011000000000000111100000000;
    wire [5:0] lut_2101_select = {
                             in_data[685],
                             in_data[157],
                             in_data[353],
                             in_data[348],
                             in_data[238],
                             in_data[26]};
    
    wire lut_2101_out = lut_2101_table[lut_2101_select];
    
    generate
    if ( USE_REG ) begin : ff_2101
        reg   lut_2101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2101_ff <= lut_2101_out;
            end
        end
        
        assign out_data[2101] = lut_2101_ff;
    end
    else begin : no_ff_2101
        assign out_data[2101] = lut_2101_out;
    end
    endgenerate
    
    
    
    // LUT : 2102
    wire [63:0] lut_2102_table = 64'b1111111111111111111111111111111111111101011111000001000001110000;
    wire [5:0] lut_2102_select = {
                             in_data[568],
                             in_data[95],
                             in_data[389],
                             in_data[160],
                             in_data[180],
                             in_data[741]};
    
    wire lut_2102_out = lut_2102_table[lut_2102_select];
    
    generate
    if ( USE_REG ) begin : ff_2102
        reg   lut_2102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2102_ff <= lut_2102_out;
            end
        end
        
        assign out_data[2102] = lut_2102_ff;
    end
    else begin : no_ff_2102
        assign out_data[2102] = lut_2102_out;
    end
    endgenerate
    
    
    
    // LUT : 2103
    wire [63:0] lut_2103_table = 64'b1010101000000000101010100000000010101010000010101010101000001010;
    wire [5:0] lut_2103_select = {
                             in_data[484],
                             in_data[3],
                             in_data[381],
                             in_data[190],
                             in_data[765],
                             in_data[183]};
    
    wire lut_2103_out = lut_2103_table[lut_2103_select];
    
    generate
    if ( USE_REG ) begin : ff_2103
        reg   lut_2103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2103_ff <= lut_2103_out;
            end
        end
        
        assign out_data[2103] = lut_2103_ff;
    end
    else begin : no_ff_2103
        assign out_data[2103] = lut_2103_out;
    end
    endgenerate
    
    
    
    // LUT : 2104
    wire [63:0] lut_2104_table = 64'b1111111111111100111111111111110011111100111100001111110011111000;
    wire [5:0] lut_2104_select = {
                             in_data[570],
                             in_data[450],
                             in_data[68],
                             in_data[540],
                             in_data[656],
                             in_data[47]};
    
    wire lut_2104_out = lut_2104_table[lut_2104_select];
    
    generate
    if ( USE_REG ) begin : ff_2104
        reg   lut_2104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2104_ff <= lut_2104_out;
            end
        end
        
        assign out_data[2104] = lut_2104_ff;
    end
    else begin : no_ff_2104
        assign out_data[2104] = lut_2104_out;
    end
    endgenerate
    
    
    
    // LUT : 2105
    wire [63:0] lut_2105_table = 64'b1111010101010001111111111101000011110101010100011111111111110000;
    wire [5:0] lut_2105_select = {
                             in_data[309],
                             in_data[159],
                             in_data[184],
                             in_data[121],
                             in_data[588],
                             in_data[518]};
    
    wire lut_2105_out = lut_2105_table[lut_2105_select];
    
    generate
    if ( USE_REG ) begin : ff_2105
        reg   lut_2105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2105_ff <= lut_2105_out;
            end
        end
        
        assign out_data[2105] = lut_2105_ff;
    end
    else begin : no_ff_2105
        assign out_data[2105] = lut_2105_out;
    end
    endgenerate
    
    
    
    // LUT : 2106
    wire [63:0] lut_2106_table = 64'b0000000000000000010101010000000011111111000000001111111100000000;
    wire [5:0] lut_2106_select = {
                             in_data[323],
                             in_data[608],
                             in_data[158],
                             in_data[254],
                             in_data[641],
                             in_data[452]};
    
    wire lut_2106_out = lut_2106_table[lut_2106_select];
    
    generate
    if ( USE_REG ) begin : ff_2106
        reg   lut_2106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2106_ff <= lut_2106_out;
            end
        end
        
        assign out_data[2106] = lut_2106_ff;
    end
    else begin : no_ff_2106
        assign out_data[2106] = lut_2106_out;
    end
    endgenerate
    
    
    
    // LUT : 2107
    wire [63:0] lut_2107_table = 64'b1010111110101111100011111010111100001110000011100000100000000000;
    wire [5:0] lut_2107_select = {
                             in_data[440],
                             in_data[163],
                             in_data[767],
                             in_data[73],
                             in_data[732],
                             in_data[455]};
    
    wire lut_2107_out = lut_2107_table[lut_2107_select];
    
    generate
    if ( USE_REG ) begin : ff_2107
        reg   lut_2107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2107_ff <= lut_2107_out;
            end
        end
        
        assign out_data[2107] = lut_2107_ff;
    end
    else begin : no_ff_2107
        assign out_data[2107] = lut_2107_out;
    end
    endgenerate
    
    
    
    // LUT : 2108
    wire [63:0] lut_2108_table = 64'b1010101011101110111111111111111111101100111011101100111011001111;
    wire [5:0] lut_2108_select = {
                             in_data[344],
                             in_data[627],
                             in_data[639],
                             in_data[120],
                             in_data[341],
                             in_data[331]};
    
    wire lut_2108_out = lut_2108_table[lut_2108_select];
    
    generate
    if ( USE_REG ) begin : ff_2108
        reg   lut_2108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2108_ff <= lut_2108_out;
            end
        end
        
        assign out_data[2108] = lut_2108_ff;
    end
    else begin : no_ff_2108
        assign out_data[2108] = lut_2108_out;
    end
    endgenerate
    
    
    
    // LUT : 2109
    wire [63:0] lut_2109_table = 64'b1111111111111111110011001100110011111111111111111100110011001100;
    wire [5:0] lut_2109_select = {
                             in_data[702],
                             in_data[385],
                             in_data[266],
                             in_data[477],
                             in_data[637],
                             in_data[114]};
    
    wire lut_2109_out = lut_2109_table[lut_2109_select];
    
    generate
    if ( USE_REG ) begin : ff_2109
        reg   lut_2109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2109_ff <= lut_2109_out;
            end
        end
        
        assign out_data[2109] = lut_2109_ff;
    end
    else begin : no_ff_2109
        assign out_data[2109] = lut_2109_out;
    end
    endgenerate
    
    
    
    // LUT : 2110
    wire [63:0] lut_2110_table = 64'b1111010100000000111101110000000011110101000000001111010100000000;
    wire [5:0] lut_2110_select = {
                             in_data[728],
                             in_data[5],
                             in_data[461],
                             in_data[447],
                             in_data[779],
                             in_data[691]};
    
    wire lut_2110_out = lut_2110_table[lut_2110_select];
    
    generate
    if ( USE_REG ) begin : ff_2110
        reg   lut_2110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2110_ff <= lut_2110_out;
            end
        end
        
        assign out_data[2110] = lut_2110_ff;
    end
    else begin : no_ff_2110
        assign out_data[2110] = lut_2110_out;
    end
    endgenerate
    
    
    
    // LUT : 2111
    wire [63:0] lut_2111_table = 64'b0000000000000000000100000000000000000000000000000011111100001111;
    wire [5:0] lut_2111_select = {
                             in_data[522],
                             in_data[386],
                             in_data[352],
                             in_data[374],
                             in_data[507],
                             in_data[587]};
    
    wire lut_2111_out = lut_2111_table[lut_2111_select];
    
    generate
    if ( USE_REG ) begin : ff_2111
        reg   lut_2111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2111_ff <= lut_2111_out;
            end
        end
        
        assign out_data[2111] = lut_2111_ff;
    end
    else begin : no_ff_2111
        assign out_data[2111] = lut_2111_out;
    end
    endgenerate
    
    
    
    // LUT : 2112
    wire [63:0] lut_2112_table = 64'b1111110011111100111111111111111111111100111111001111110011111111;
    wire [5:0] lut_2112_select = {
                             in_data[501],
                             in_data[299],
                             in_data[57],
                             in_data[630],
                             in_data[277],
                             in_data[88]};
    
    wire lut_2112_out = lut_2112_table[lut_2112_select];
    
    generate
    if ( USE_REG ) begin : ff_2112
        reg   lut_2112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2112_ff <= lut_2112_out;
            end
        end
        
        assign out_data[2112] = lut_2112_ff;
    end
    else begin : no_ff_2112
        assign out_data[2112] = lut_2112_out;
    end
    endgenerate
    
    
    
    // LUT : 2113
    wire [63:0] lut_2113_table = 64'b1110111011101110111011101110111011101110111011101110111011101110;
    wire [5:0] lut_2113_select = {
                             in_data[165],
                             in_data[125],
                             in_data[116],
                             in_data[94],
                             in_data[319],
                             in_data[97]};
    
    wire lut_2113_out = lut_2113_table[lut_2113_select];
    
    generate
    if ( USE_REG ) begin : ff_2113
        reg   lut_2113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2113_ff <= lut_2113_out;
            end
        end
        
        assign out_data[2113] = lut_2113_ff;
    end
    else begin : no_ff_2113
        assign out_data[2113] = lut_2113_out;
    end
    endgenerate
    
    
    
    // LUT : 2114
    wire [63:0] lut_2114_table = 64'b1011101111111111001000101011101111111111111111110010001010101010;
    wire [5:0] lut_2114_select = {
                             in_data[380],
                             in_data[653],
                             in_data[276],
                             in_data[17],
                             in_data[715],
                             in_data[709]};
    
    wire lut_2114_out = lut_2114_table[lut_2114_select];
    
    generate
    if ( USE_REG ) begin : ff_2114
        reg   lut_2114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2114_ff <= lut_2114_out;
            end
        end
        
        assign out_data[2114] = lut_2114_ff;
    end
    else begin : no_ff_2114
        assign out_data[2114] = lut_2114_out;
    end
    endgenerate
    
    
    
    // LUT : 2115
    wire [63:0] lut_2115_table = 64'b0000000000000000000000000000000000000000000000000000111100001111;
    wire [5:0] lut_2115_select = {
                             in_data[186],
                             in_data[622],
                             in_data[419],
                             in_data[594],
                             in_data[167],
                             in_data[393]};
    
    wire lut_2115_out = lut_2115_table[lut_2115_select];
    
    generate
    if ( USE_REG ) begin : ff_2115
        reg   lut_2115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2115_ff <= lut_2115_out;
            end
        end
        
        assign out_data[2115] = lut_2115_ff;
    end
    else begin : no_ff_2115
        assign out_data[2115] = lut_2115_out;
    end
    endgenerate
    
    
    
    // LUT : 2116
    wire [63:0] lut_2116_table = 64'b1111111111111111010000001111111111111111111111110100000011111111;
    wire [5:0] lut_2116_select = {
                             in_data[640],
                             in_data[684],
                             in_data[324],
                             in_data[103],
                             in_data[438],
                             in_data[689]};
    
    wire lut_2116_out = lut_2116_table[lut_2116_select];
    
    generate
    if ( USE_REG ) begin : ff_2116
        reg   lut_2116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2116_ff <= lut_2116_out;
            end
        end
        
        assign out_data[2116] = lut_2116_ff;
    end
    else begin : no_ff_2116
        assign out_data[2116] = lut_2116_out;
    end
    endgenerate
    
    
    
    // LUT : 2117
    wire [63:0] lut_2117_table = 64'b1111111111011101110111011100110011001100010011000100010001000100;
    wire [5:0] lut_2117_select = {
                             in_data[628],
                             in_data[231],
                             in_data[638],
                             in_data[111],
                             in_data[572],
                             in_data[619]};
    
    wire lut_2117_out = lut_2117_table[lut_2117_select];
    
    generate
    if ( USE_REG ) begin : ff_2117
        reg   lut_2117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2117_ff <= lut_2117_out;
            end
        end
        
        assign out_data[2117] = lut_2117_ff;
    end
    else begin : no_ff_2117
        assign out_data[2117] = lut_2117_out;
    end
    endgenerate
    
    
    
    // LUT : 2118
    wire [63:0] lut_2118_table = 64'b1110110011111111111011001111111111101100111111111110110011111111;
    wire [5:0] lut_2118_select = {
                             in_data[308],
                             in_data[11],
                             in_data[545],
                             in_data[668],
                             in_data[304],
                             in_data[771]};
    
    wire lut_2118_out = lut_2118_table[lut_2118_select];
    
    generate
    if ( USE_REG ) begin : ff_2118
        reg   lut_2118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2118_ff <= lut_2118_out;
            end
        end
        
        assign out_data[2118] = lut_2118_ff;
    end
    else begin : no_ff_2118
        assign out_data[2118] = lut_2118_out;
    end
    endgenerate
    
    
    
    // LUT : 2119
    wire [63:0] lut_2119_table = 64'b0000000000000000001100110000000000000000000000001111111111001111;
    wire [5:0] lut_2119_select = {
                             in_data[291],
                             in_data[661],
                             in_data[327],
                             in_data[75],
                             in_data[124],
                             in_data[335]};
    
    wire lut_2119_out = lut_2119_table[lut_2119_select];
    
    generate
    if ( USE_REG ) begin : ff_2119
        reg   lut_2119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2119_ff <= lut_2119_out;
            end
        end
        
        assign out_data[2119] = lut_2119_ff;
    end
    else begin : no_ff_2119
        assign out_data[2119] = lut_2119_out;
    end
    endgenerate
    
    
    
    // LUT : 2120
    wire [63:0] lut_2120_table = 64'b1111111100001100111111110000110011111111000011001110111100001100;
    wire [5:0] lut_2120_select = {
                             in_data[711],
                             in_data[647],
                             in_data[325],
                             in_data[625],
                             in_data[473],
                             in_data[9]};
    
    wire lut_2120_out = lut_2120_table[lut_2120_select];
    
    generate
    if ( USE_REG ) begin : ff_2120
        reg   lut_2120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2120_ff <= lut_2120_out;
            end
        end
        
        assign out_data[2120] = lut_2120_ff;
    end
    else begin : no_ff_2120
        assign out_data[2120] = lut_2120_out;
    end
    endgenerate
    
    
    
    // LUT : 2121
    wire [63:0] lut_2121_table = 64'b1111111111111111000000000000101011111111111111110000000000000000;
    wire [5:0] lut_2121_select = {
                             in_data[757],
                             in_data[467],
                             in_data[227],
                             in_data[214],
                             in_data[337],
                             in_data[228]};
    
    wire lut_2121_out = lut_2121_table[lut_2121_select];
    
    generate
    if ( USE_REG ) begin : ff_2121
        reg   lut_2121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2121_ff <= lut_2121_out;
            end
        end
        
        assign out_data[2121] = lut_2121_ff;
    end
    else begin : no_ff_2121
        assign out_data[2121] = lut_2121_out;
    end
    endgenerate
    
    
    
    // LUT : 2122
    wire [63:0] lut_2122_table = 64'b1010101010101010101010101010101010100010001000101010001010100010;
    wire [5:0] lut_2122_select = {
                             in_data[706],
                             in_data[615],
                             in_data[90],
                             in_data[504],
                             in_data[286],
                             in_data[411]};
    
    wire lut_2122_out = lut_2122_table[lut_2122_select];
    
    generate
    if ( USE_REG ) begin : ff_2122
        reg   lut_2122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2122_ff <= lut_2122_out;
            end
        end
        
        assign out_data[2122] = lut_2122_ff;
    end
    else begin : no_ff_2122
        assign out_data[2122] = lut_2122_out;
    end
    endgenerate
    
    
    
    // LUT : 2123
    wire [63:0] lut_2123_table = 64'b0000111000000000000011110000010000001111000000000101111100000100;
    wire [5:0] lut_2123_select = {
                             in_data[232],
                             in_data[396],
                             in_data[377],
                             in_data[525],
                             in_data[609],
                             in_data[553]};
    
    wire lut_2123_out = lut_2123_table[lut_2123_select];
    
    generate
    if ( USE_REG ) begin : ff_2123
        reg   lut_2123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2123_ff <= lut_2123_out;
            end
        end
        
        assign out_data[2123] = lut_2123_ff;
    end
    else begin : no_ff_2123
        assign out_data[2123] = lut_2123_out;
    end
    endgenerate
    
    
    
    // LUT : 2124
    wire [63:0] lut_2124_table = 64'b1111111111111111111111111111111101011101010111010101110101010101;
    wire [5:0] lut_2124_select = {
                             in_data[708],
                             in_data[763],
                             in_data[23],
                             in_data[223],
                             in_data[118],
                             in_data[626]};
    
    wire lut_2124_out = lut_2124_table[lut_2124_select];
    
    generate
    if ( USE_REG ) begin : ff_2124
        reg   lut_2124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2124_ff <= lut_2124_out;
            end
        end
        
        assign out_data[2124] = lut_2124_ff;
    end
    else begin : no_ff_2124
        assign out_data[2124] = lut_2124_out;
    end
    endgenerate
    
    
    
    // LUT : 2125
    wire [63:0] lut_2125_table = 64'b1111111111111111000011010000010111111111000011110000010100000000;
    wire [5:0] lut_2125_select = {
                             in_data[735],
                             in_data[521],
                             in_data[480],
                             in_data[427],
                             in_data[56],
                             in_data[274]};
    
    wire lut_2125_out = lut_2125_table[lut_2125_select];
    
    generate
    if ( USE_REG ) begin : ff_2125
        reg   lut_2125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2125_ff <= lut_2125_out;
            end
        end
        
        assign out_data[2125] = lut_2125_ff;
    end
    else begin : no_ff_2125
        assign out_data[2125] = lut_2125_out;
    end
    endgenerate
    
    
    
    // LUT : 2126
    wire [63:0] lut_2126_table = 64'b1111111111111111111111111111111110100000101000001010000010100000;
    wire [5:0] lut_2126_select = {
                             in_data[548],
                             in_data[783],
                             in_data[643],
                             in_data[300],
                             in_data[750],
                             in_data[93]};
    
    wire lut_2126_out = lut_2126_table[lut_2126_select];
    
    generate
    if ( USE_REG ) begin : ff_2126
        reg   lut_2126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2126_ff <= lut_2126_out;
            end
        end
        
        assign out_data[2126] = lut_2126_ff;
    end
    else begin : no_ff_2126
        assign out_data[2126] = lut_2126_out;
    end
    endgenerate
    
    
    
    // LUT : 2127
    wire [63:0] lut_2127_table = 64'b0000110011111111000011001111111100000000111111000001000011111111;
    wire [5:0] lut_2127_select = {
                             in_data[482],
                             in_data[112],
                             in_data[544],
                             in_data[376],
                             in_data[314],
                             in_data[48]};
    
    wire lut_2127_out = lut_2127_table[lut_2127_select];
    
    generate
    if ( USE_REG ) begin : ff_2127
        reg   lut_2127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2127_ff <= lut_2127_out;
            end
        end
        
        assign out_data[2127] = lut_2127_ff;
    end
    else begin : no_ff_2127
        assign out_data[2127] = lut_2127_out;
    end
    endgenerate
    
    
    
    // LUT : 2128
    wire [63:0] lut_2128_table = 64'b1111111111111111111111111111111100000000000000000101010000000000;
    wire [5:0] lut_2128_select = {
                             in_data[209],
                             in_data[659],
                             in_data[508],
                             in_data[55],
                             in_data[85],
                             in_data[692]};
    
    wire lut_2128_out = lut_2128_table[lut_2128_select];
    
    generate
    if ( USE_REG ) begin : ff_2128
        reg   lut_2128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2128_ff <= lut_2128_out;
            end
        end
        
        assign out_data[2128] = lut_2128_ff;
    end
    else begin : no_ff_2128
        assign out_data[2128] = lut_2128_out;
    end
    endgenerate
    
    
    
    // LUT : 2129
    wire [63:0] lut_2129_table = 64'b1111101011110000111100001111000011110000111101011111000011110101;
    wire [5:0] lut_2129_select = {
                             in_data[511],
                             in_data[646],
                             in_data[486],
                             in_data[597],
                             in_data[169],
                             in_data[349]};
    
    wire lut_2129_out = lut_2129_table[lut_2129_select];
    
    generate
    if ( USE_REG ) begin : ff_2129
        reg   lut_2129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2129_ff <= lut_2129_out;
            end
        end
        
        assign out_data[2129] = lut_2129_ff;
    end
    else begin : no_ff_2129
        assign out_data[2129] = lut_2129_out;
    end
    endgenerate
    
    
    
    // LUT : 2130
    wire [63:0] lut_2130_table = 64'b1111111111111111000001010000000100000101000001010000010100000101;
    wire [5:0] lut_2130_select = {
                             in_data[148],
                             in_data[574],
                             in_data[394],
                             in_data[464],
                             in_data[729],
                             in_data[357]};
    
    wire lut_2130_out = lut_2130_table[lut_2130_select];
    
    generate
    if ( USE_REG ) begin : ff_2130
        reg   lut_2130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2130_ff <= lut_2130_out;
            end
        end
        
        assign out_data[2130] = lut_2130_ff;
    end
    else begin : no_ff_2130
        assign out_data[2130] = lut_2130_out;
    end
    endgenerate
    
    
    
    // LUT : 2131
    wire [63:0] lut_2131_table = 64'b0011111100111111000011110000111100111111101111110000111000001111;
    wire [5:0] lut_2131_select = {
                             in_data[773],
                             in_data[128],
                             in_data[83],
                             in_data[409],
                             in_data[485],
                             in_data[44]};
    
    wire lut_2131_out = lut_2131_table[lut_2131_select];
    
    generate
    if ( USE_REG ) begin : ff_2131
        reg   lut_2131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2131_ff <= lut_2131_out;
            end
        end
        
        assign out_data[2131] = lut_2131_ff;
    end
    else begin : no_ff_2131
        assign out_data[2131] = lut_2131_out;
    end
    endgenerate
    
    
    
    // LUT : 2132
    wire [63:0] lut_2132_table = 64'b0011001100110011001000100010001000110011001100111011101010101010;
    wire [5:0] lut_2132_select = {
                             in_data[310],
                             in_data[262],
                             in_data[307],
                             in_data[704],
                             in_data[442],
                             in_data[178]};
    
    wire lut_2132_out = lut_2132_table[lut_2132_select];
    
    generate
    if ( USE_REG ) begin : ff_2132
        reg   lut_2132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2132_ff <= lut_2132_out;
            end
        end
        
        assign out_data[2132] = lut_2132_ff;
    end
    else begin : no_ff_2132
        assign out_data[2132] = lut_2132_out;
    end
    endgenerate
    
    
    
    // LUT : 2133
    wire [63:0] lut_2133_table = 64'b0000000000000000000000000000000011011101110011001101110111001100;
    wire [5:0] lut_2133_select = {
                             in_data[707],
                             in_data[644],
                             in_data[360],
                             in_data[418],
                             in_data[298],
                             in_data[368]};
    
    wire lut_2133_out = lut_2133_table[lut_2133_select];
    
    generate
    if ( USE_REG ) begin : ff_2133
        reg   lut_2133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2133_ff <= lut_2133_out;
            end
        end
        
        assign out_data[2133] = lut_2133_ff;
    end
    else begin : no_ff_2133
        assign out_data[2133] = lut_2133_out;
    end
    endgenerate
    
    
    
    // LUT : 2134
    wire [63:0] lut_2134_table = 64'b1111111111001100110111011100110011111111110011011100110011001100;
    wire [5:0] lut_2134_select = {
                             in_data[144],
                             in_data[242],
                             in_data[220],
                             in_data[249],
                             in_data[539],
                             in_data[197]};
    
    wire lut_2134_out = lut_2134_table[lut_2134_select];
    
    generate
    if ( USE_REG ) begin : ff_2134
        reg   lut_2134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2134_ff <= lut_2134_out;
            end
        end
        
        assign out_data[2134] = lut_2134_ff;
    end
    else begin : no_ff_2134
        assign out_data[2134] = lut_2134_out;
    end
    endgenerate
    
    
    
    // LUT : 2135
    wire [63:0] lut_2135_table = 64'b0000010101011101010101011101110100000000010001000000000001000101;
    wire [5:0] lut_2135_select = {
                             in_data[526],
                             in_data[226],
                             in_data[270],
                             in_data[200],
                             in_data[569],
                             in_data[229]};
    
    wire lut_2135_out = lut_2135_table[lut_2135_select];
    
    generate
    if ( USE_REG ) begin : ff_2135
        reg   lut_2135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2135_ff <= lut_2135_out;
            end
        end
        
        assign out_data[2135] = lut_2135_ff;
    end
    else begin : no_ff_2135
        assign out_data[2135] = lut_2135_out;
    end
    endgenerate
    
    
    
    // LUT : 2136
    wire [63:0] lut_2136_table = 64'b0000000011111111000000001111111100000000111111010000000011111101;
    wire [5:0] lut_2136_select = {
                             in_data[496],
                             in_data[12],
                             in_data[289],
                             in_data[523],
                             in_data[654],
                             in_data[104]};
    
    wire lut_2136_out = lut_2136_table[lut_2136_select];
    
    generate
    if ( USE_REG ) begin : ff_2136
        reg   lut_2136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2136_ff <= lut_2136_out;
            end
        end
        
        assign out_data[2136] = lut_2136_ff;
    end
    else begin : no_ff_2136
        assign out_data[2136] = lut_2136_out;
    end
    endgenerate
    
    
    
    // LUT : 2137
    wire [63:0] lut_2137_table = 64'b0000000000110011000000000000000000110011001100110000000000110011;
    wire [5:0] lut_2137_select = {
                             in_data[551],
                             in_data[736],
                             in_data[155],
                             in_data[338],
                             in_data[610],
                             in_data[84]};
    
    wire lut_2137_out = lut_2137_table[lut_2137_select];
    
    generate
    if ( USE_REG ) begin : ff_2137
        reg   lut_2137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2137_ff <= lut_2137_out;
            end
        end
        
        assign out_data[2137] = lut_2137_ff;
    end
    else begin : no_ff_2137
        assign out_data[2137] = lut_2137_out;
    end
    endgenerate
    
    
    
    // LUT : 2138
    wire [63:0] lut_2138_table = 64'b1111111101110101111111110111111101010101010101010101010101010101;
    wire [5:0] lut_2138_select = {
                             in_data[175],
                             in_data[34],
                             in_data[251],
                             in_data[1],
                             in_data[59],
                             in_data[462]};
    
    wire lut_2138_out = lut_2138_table[lut_2138_select];
    
    generate
    if ( USE_REG ) begin : ff_2138
        reg   lut_2138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2138_ff <= lut_2138_out;
            end
        end
        
        assign out_data[2138] = lut_2138_ff;
    end
    else begin : no_ff_2138
        assign out_data[2138] = lut_2138_out;
    end
    endgenerate
    
    
    
    // LUT : 2139
    wire [63:0] lut_2139_table = 64'b1111111111110010111111111111001111111111101000001111111110110000;
    wire [5:0] lut_2139_select = {
                             in_data[426],
                             in_data[290],
                             in_data[481],
                             in_data[575],
                             in_data[361],
                             in_data[96]};
    
    wire lut_2139_out = lut_2139_table[lut_2139_select];
    
    generate
    if ( USE_REG ) begin : ff_2139
        reg   lut_2139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2139_ff <= lut_2139_out;
            end
        end
        
        assign out_data[2139] = lut_2139_ff;
    end
    else begin : no_ff_2139
        assign out_data[2139] = lut_2139_out;
    end
    endgenerate
    
    
    
    // LUT : 2140
    wire [63:0] lut_2140_table = 64'b0001001100110011001000010011001100000000111100110000000011110011;
    wire [5:0] lut_2140_select = {
                             in_data[211],
                             in_data[43],
                             in_data[132],
                             in_data[383],
                             in_data[541],
                             in_data[751]};
    
    wire lut_2140_out = lut_2140_table[lut_2140_select];
    
    generate
    if ( USE_REG ) begin : ff_2140
        reg   lut_2140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2140_ff <= lut_2140_out;
            end
        end
        
        assign out_data[2140] = lut_2140_ff;
    end
    else begin : no_ff_2140
        assign out_data[2140] = lut_2140_out;
    end
    endgenerate
    
    
    
    // LUT : 2141
    wire [63:0] lut_2141_table = 64'b0011001100110011001100110011011100010001001100110000000000010001;
    wire [5:0] lut_2141_select = {
                             in_data[660],
                             in_data[230],
                             in_data[676],
                             in_data[505],
                             in_data[265],
                             in_data[137]};
    
    wire lut_2141_out = lut_2141_table[lut_2141_select];
    
    generate
    if ( USE_REG ) begin : ff_2141
        reg   lut_2141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2141_ff <= lut_2141_out;
            end
        end
        
        assign out_data[2141] = lut_2141_ff;
    end
    else begin : no_ff_2141
        assign out_data[2141] = lut_2141_out;
    end
    endgenerate
    
    
    
    // LUT : 2142
    wire [63:0] lut_2142_table = 64'b1111000011110101111101011111010111110000111100001111000011110000;
    wire [5:0] lut_2142_select = {
                             in_data[405],
                             in_data[726],
                             in_data[421],
                             in_data[469],
                             in_data[224],
                             in_data[744]};
    
    wire lut_2142_out = lut_2142_table[lut_2142_select];
    
    generate
    if ( USE_REG ) begin : ff_2142
        reg   lut_2142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2142_ff <= lut_2142_out;
            end
        end
        
        assign out_data[2142] = lut_2142_ff;
    end
    else begin : no_ff_2142
        assign out_data[2142] = lut_2142_out;
    end
    endgenerate
    
    
    
    // LUT : 2143
    wire [63:0] lut_2143_table = 64'b0001000100010001000000000001000011001100110011001100110011001100;
    wire [5:0] lut_2143_select = {
                             in_data[537],
                             in_data[694],
                             in_data[422],
                             in_data[696],
                             in_data[517],
                             in_data[451]};
    
    wire lut_2143_out = lut_2143_table[lut_2143_select];
    
    generate
    if ( USE_REG ) begin : ff_2143
        reg   lut_2143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2143_ff <= lut_2143_out;
            end
        end
        
        assign out_data[2143] = lut_2143_ff;
    end
    else begin : no_ff_2143
        assign out_data[2143] = lut_2143_out;
    end
    endgenerate
    
    
    
    // LUT : 2144
    wire [63:0] lut_2144_table = 64'b0000000011111111000000001111111100000000111111110000000011111111;
    wire [5:0] lut_2144_select = {
                             in_data[710],
                             in_data[693],
                             in_data[268],
                             in_data[761],
                             in_data[586],
                             in_data[69]};
    
    wire lut_2144_out = lut_2144_table[lut_2144_select];
    
    generate
    if ( USE_REG ) begin : ff_2144
        reg   lut_2144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2144_ff <= lut_2144_out;
            end
        end
        
        assign out_data[2144] = lut_2144_ff;
    end
    else begin : no_ff_2144
        assign out_data[2144] = lut_2144_out;
    end
    endgenerate
    
    
    
    // LUT : 2145
    wire [63:0] lut_2145_table = 64'b1111111111111111111111111111111111111111111111110000110000001100;
    wire [5:0] lut_2145_select = {
                             in_data[416],
                             in_data[187],
                             in_data[478],
                             in_data[687],
                             in_data[201],
                             in_data[102]};
    
    wire lut_2145_out = lut_2145_table[lut_2145_select];
    
    generate
    if ( USE_REG ) begin : ff_2145
        reg   lut_2145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2145_ff <= lut_2145_out;
            end
        end
        
        assign out_data[2145] = lut_2145_ff;
    end
    else begin : no_ff_2145
        assign out_data[2145] = lut_2145_out;
    end
    endgenerate
    
    
    
    // LUT : 2146
    wire [63:0] lut_2146_table = 64'b0101010111010101010101011101110011010101110101010101010111011100;
    wire [5:0] lut_2146_select = {
                             in_data[560],
                             in_data[493],
                             in_data[494],
                             in_data[436],
                             in_data[333],
                             in_data[375]};
    
    wire lut_2146_out = lut_2146_table[lut_2146_select];
    
    generate
    if ( USE_REG ) begin : ff_2146
        reg   lut_2146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2146_ff <= lut_2146_out;
            end
        end
        
        assign out_data[2146] = lut_2146_ff;
    end
    else begin : no_ff_2146
        assign out_data[2146] = lut_2146_out;
    end
    endgenerate
    
    
    
    // LUT : 2147
    wire [63:0] lut_2147_table = 64'b1010000010100000101000001010000011110101111101011111010111110101;
    wire [5:0] lut_2147_select = {
                             in_data[402],
                             in_data[62],
                             in_data[697],
                             in_data[205],
                             in_data[115],
                             in_data[635]};
    
    wire lut_2147_out = lut_2147_table[lut_2147_select];
    
    generate
    if ( USE_REG ) begin : ff_2147
        reg   lut_2147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2147_ff <= lut_2147_out;
            end
        end
        
        assign out_data[2147] = lut_2147_ff;
    end
    else begin : no_ff_2147
        assign out_data[2147] = lut_2147_out;
    end
    endgenerate
    
    
    
    // LUT : 2148
    wire [63:0] lut_2148_table = 64'b1111111111111111111111111111111111101111101011111010111110101111;
    wire [5:0] lut_2148_select = {
                             in_data[74],
                             in_data[279],
                             in_data[89],
                             in_data[240],
                             in_data[764],
                             in_data[202]};
    
    wire lut_2148_out = lut_2148_table[lut_2148_select];
    
    generate
    if ( USE_REG ) begin : ff_2148
        reg   lut_2148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2148_ff <= lut_2148_out;
            end
        end
        
        assign out_data[2148] = lut_2148_ff;
    end
    else begin : no_ff_2148
        assign out_data[2148] = lut_2148_out;
    end
    endgenerate
    
    
    
    // LUT : 2149
    wire [63:0] lut_2149_table = 64'b0001000101111111000000000000000000010001011111110000000000000000;
    wire [5:0] lut_2149_select = {
                             in_data[81],
                             in_data[126],
                             in_data[680],
                             in_data[770],
                             in_data[234],
                             in_data[679]};
    
    wire lut_2149_out = lut_2149_table[lut_2149_select];
    
    generate
    if ( USE_REG ) begin : ff_2149
        reg   lut_2149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2149_ff <= lut_2149_out;
            end
        end
        
        assign out_data[2149] = lut_2149_ff;
    end
    else begin : no_ff_2149
        assign out_data[2149] = lut_2149_out;
    end
    endgenerate
    
    
    
    // LUT : 2150
    wire [63:0] lut_2150_table = 64'b0100000001000000010111000101110001001100010011001101111111011111;
    wire [5:0] lut_2150_select = {
                             in_data[435],
                             in_data[743],
                             in_data[51],
                             in_data[192],
                             in_data[500],
                             in_data[216]};
    
    wire lut_2150_out = lut_2150_table[lut_2150_select];
    
    generate
    if ( USE_REG ) begin : ff_2150
        reg   lut_2150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2150_ff <= lut_2150_out;
            end
        end
        
        assign out_data[2150] = lut_2150_ff;
    end
    else begin : no_ff_2150
        assign out_data[2150] = lut_2150_out;
    end
    endgenerate
    
    
    
    // LUT : 2151
    wire [63:0] lut_2151_table = 64'b1010101010111111000000000010101110101010101111110000000010101010;
    wire [5:0] lut_2151_select = {
                             in_data[58],
                             in_data[78],
                             in_data[747],
                             in_data[37],
                             in_data[558],
                             in_data[106]};
    
    wire lut_2151_out = lut_2151_table[lut_2151_select];
    
    generate
    if ( USE_REG ) begin : ff_2151
        reg   lut_2151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2151_ff <= lut_2151_out;
            end
        end
        
        assign out_data[2151] = lut_2151_ff;
    end
    else begin : no_ff_2151
        assign out_data[2151] = lut_2151_out;
    end
    endgenerate
    
    
    
    // LUT : 2152
    wire [63:0] lut_2152_table = 64'b1111101011111010111110101111101010111010111110101010101011111010;
    wire [5:0] lut_2152_select = {
                             in_data[671],
                             in_data[52],
                             in_data[470],
                             in_data[194],
                             in_data[225],
                             in_data[550]};
    
    wire lut_2152_out = lut_2152_table[lut_2152_select];
    
    generate
    if ( USE_REG ) begin : ff_2152
        reg   lut_2152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2152_ff <= lut_2152_out;
            end
        end
        
        assign out_data[2152] = lut_2152_ff;
    end
    else begin : no_ff_2152
        assign out_data[2152] = lut_2152_out;
    end
    endgenerate
    
    
    
    // LUT : 2153
    wire [63:0] lut_2153_table = 64'b0100111111001110010011011100111001001111010011110100111101001111;
    wire [5:0] lut_2153_select = {
                             in_data[358],
                             in_data[590],
                             in_data[152],
                             in_data[317],
                             in_data[218],
                             in_data[176]};
    
    wire lut_2153_out = lut_2153_table[lut_2153_select];
    
    generate
    if ( USE_REG ) begin : ff_2153
        reg   lut_2153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2153_ff <= lut_2153_out;
            end
        end
        
        assign out_data[2153] = lut_2153_ff;
    end
    else begin : no_ff_2153
        assign out_data[2153] = lut_2153_out;
    end
    endgenerate
    
    
    
    // LUT : 2154
    wire [63:0] lut_2154_table = 64'b0000000000001111000000000000111111111111111111111100111111111111;
    wire [5:0] lut_2154_select = {
                             in_data[297],
                             in_data[14],
                             in_data[549],
                             in_data[600],
                             in_data[133],
                             in_data[33]};
    
    wire lut_2154_out = lut_2154_table[lut_2154_select];
    
    generate
    if ( USE_REG ) begin : ff_2154
        reg   lut_2154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2154_ff <= lut_2154_out;
            end
        end
        
        assign out_data[2154] = lut_2154_ff;
    end
    else begin : no_ff_2154
        assign out_data[2154] = lut_2154_out;
    end
    endgenerate
    
    
    
    // LUT : 2155
    wire [63:0] lut_2155_table = 64'b1000100000000000101010100000000011101110101010101111111110101010;
    wire [5:0] lut_2155_select = {
                             in_data[566],
                             in_data[311],
                             in_data[305],
                             in_data[278],
                             in_data[92],
                             in_data[492]};
    
    wire lut_2155_out = lut_2155_table[lut_2155_select];
    
    generate
    if ( USE_REG ) begin : ff_2155
        reg   lut_2155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2155_ff <= lut_2155_out;
            end
        end
        
        assign out_data[2155] = lut_2155_ff;
    end
    else begin : no_ff_2155
        assign out_data[2155] = lut_2155_out;
    end
    endgenerate
    
    
    
    // LUT : 2156
    wire [63:0] lut_2156_table = 64'b0000000000000000001010101010111000000000000000000000111100001111;
    wire [5:0] lut_2156_select = {
                             in_data[293],
                             in_data[245],
                             in_data[674],
                             in_data[127],
                             in_data[110],
                             in_data[495]};
    
    wire lut_2156_out = lut_2156_table[lut_2156_select];
    
    generate
    if ( USE_REG ) begin : ff_2156
        reg   lut_2156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2156_ff <= lut_2156_out;
            end
        end
        
        assign out_data[2156] = lut_2156_ff;
    end
    else begin : no_ff_2156
        assign out_data[2156] = lut_2156_out;
    end
    endgenerate
    
    
    
    // LUT : 2157
    wire [63:0] lut_2157_table = 64'b1010000011111111111100001111111100000000111100000000000011110001;
    wire [5:0] lut_2157_select = {
                             in_data[564],
                             in_data[134],
                             in_data[713],
                             in_data[122],
                             in_data[19],
                             in_data[430]};
    
    wire lut_2157_out = lut_2157_table[lut_2157_select];
    
    generate
    if ( USE_REG ) begin : ff_2157
        reg   lut_2157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2157_ff <= lut_2157_out;
            end
        end
        
        assign out_data[2157] = lut_2157_ff;
    end
    else begin : no_ff_2157
        assign out_data[2157] = lut_2157_out;
    end
    endgenerate
    
    
    
    // LUT : 2158
    wire [63:0] lut_2158_table = 64'b1010101010101010101010101010101010101010101010101010101010101010;
    wire [5:0] lut_2158_select = {
                             in_data[514],
                             in_data[663],
                             in_data[22],
                             in_data[70],
                             in_data[745],
                             in_data[439]};
    
    wire lut_2158_out = lut_2158_table[lut_2158_select];
    
    generate
    if ( USE_REG ) begin : ff_2158
        reg   lut_2158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2158_ff <= lut_2158_out;
            end
        end
        
        assign out_data[2158] = lut_2158_ff;
    end
    else begin : no_ff_2158
        assign out_data[2158] = lut_2158_out;
    end
    endgenerate
    
    
    
    // LUT : 2159
    wire [63:0] lut_2159_table = 64'b1111111111011101111100011100010011111111110111011111000111000100;
    wire [5:0] lut_2159_select = {
                             in_data[63],
                             in_data[459],
                             in_data[235],
                             in_data[458],
                             in_data[179],
                             in_data[195]};
    
    wire lut_2159_out = lut_2159_table[lut_2159_select];
    
    generate
    if ( USE_REG ) begin : ff_2159
        reg   lut_2159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2159_ff <= lut_2159_out;
            end
        end
        
        assign out_data[2159] = lut_2159_ff;
    end
    else begin : no_ff_2159
        assign out_data[2159] = lut_2159_out;
    end
    endgenerate
    
    
    
    // LUT : 2160
    wire [63:0] lut_2160_table = 64'b0000100011111111000000000000110000000000111111110000000000001101;
    wire [5:0] lut_2160_select = {
                             in_data[49],
                             in_data[373],
                             in_data[634],
                             in_data[542],
                             in_data[695],
                             in_data[0]};
    
    wire lut_2160_out = lut_2160_table[lut_2160_select];
    
    generate
    if ( USE_REG ) begin : ff_2160
        reg   lut_2160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2160_ff <= lut_2160_out;
            end
        end
        
        assign out_data[2160] = lut_2160_ff;
    end
    else begin : no_ff_2160
        assign out_data[2160] = lut_2160_out;
    end
    endgenerate
    
    
    
    // LUT : 2161
    wire [63:0] lut_2161_table = 64'b1101110111001100010111010000010011011101110011000100010001000100;
    wire [5:0] lut_2161_select = {
                             in_data[399],
                             in_data[453],
                             in_data[466],
                             in_data[86],
                             in_data[414],
                             in_data[580]};
    
    wire lut_2161_out = lut_2161_table[lut_2161_select];
    
    generate
    if ( USE_REG ) begin : ff_2161
        reg   lut_2161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2161_ff <= lut_2161_out;
            end
        end
        
        assign out_data[2161] = lut_2161_ff;
    end
    else begin : no_ff_2161
        assign out_data[2161] = lut_2161_out;
    end
    endgenerate
    
    
    
    // LUT : 2162
    wire [63:0] lut_2162_table = 64'b1100110011001100111111111111111111001100110011001111111111111111;
    wire [5:0] lut_2162_select = {
                             in_data[740],
                             in_data[239],
                             in_data[166],
                             in_data[256],
                             in_data[258],
                             in_data[206]};
    
    wire lut_2162_out = lut_2162_table[lut_2162_select];
    
    generate
    if ( USE_REG ) begin : ff_2162
        reg   lut_2162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2162_ff <= lut_2162_out;
            end
        end
        
        assign out_data[2162] = lut_2162_ff;
    end
    else begin : no_ff_2162
        assign out_data[2162] = lut_2162_out;
    end
    endgenerate
    
    
    
    // LUT : 2163
    wire [63:0] lut_2163_table = 64'b0000101000001010000010100000101000001011001010110000101100001011;
    wire [5:0] lut_2163_select = {
                             in_data[718],
                             in_data[246],
                             in_data[752],
                             in_data[519],
                             in_data[204],
                             in_data[571]};
    
    wire lut_2163_out = lut_2163_table[lut_2163_select];
    
    generate
    if ( USE_REG ) begin : ff_2163
        reg   lut_2163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2163_ff <= lut_2163_out;
            end
        end
        
        assign out_data[2163] = lut_2163_ff;
    end
    else begin : no_ff_2163
        assign out_data[2163] = lut_2163_out;
    end
    endgenerate
    
    
    
    // LUT : 2164
    wire [63:0] lut_2164_table = 64'b1111111111111111111111111111111111111111111111111111101011111010;
    wire [5:0] lut_2164_select = {
                             in_data[275],
                             in_data[203],
                             in_data[145],
                             in_data[147],
                             in_data[350],
                             in_data[681]};
    
    wire lut_2164_out = lut_2164_table[lut_2164_select];
    
    generate
    if ( USE_REG ) begin : ff_2164
        reg   lut_2164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2164_ff <= lut_2164_out;
            end
        end
        
        assign out_data[2164] = lut_2164_ff;
    end
    else begin : no_ff_2164
        assign out_data[2164] = lut_2164_out;
    end
    endgenerate
    
    
    
    // LUT : 2165
    wire [63:0] lut_2165_table = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [5:0] lut_2165_select = {
                             in_data[658],
                             in_data[620],
                             in_data[28],
                             in_data[645],
                             in_data[129],
                             in_data[648]};
    
    wire lut_2165_out = lut_2165_table[lut_2165_select];
    
    generate
    if ( USE_REG ) begin : ff_2165
        reg   lut_2165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2165_ff <= lut_2165_out;
            end
        end
        
        assign out_data[2165] = lut_2165_ff;
    end
    else begin : no_ff_2165
        assign out_data[2165] = lut_2165_out;
    end
    endgenerate
    
    
    
    // LUT : 2166
    wire [63:0] lut_2166_table = 64'b1010001000110011101010101011001111101110010001001110111001110100;
    wire [5:0] lut_2166_select = {
                             in_data[384],
                             in_data[32],
                             in_data[425],
                             in_data[756],
                             in_data[287],
                             in_data[652]};
    
    wire lut_2166_out = lut_2166_table[lut_2166_select];
    
    generate
    if ( USE_REG ) begin : ff_2166
        reg   lut_2166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2166_ff <= lut_2166_out;
            end
        end
        
        assign out_data[2166] = lut_2166_ff;
    end
    else begin : no_ff_2166
        assign out_data[2166] = lut_2166_out;
    end
    endgenerate
    
    
    
    // LUT : 2167
    wire [63:0] lut_2167_table = 64'b0000000000101111000000000010111100111111000011110010111100101111;
    wire [5:0] lut_2167_select = {
                             in_data[215],
                             in_data[198],
                             in_data[408],
                             in_data[579],
                             in_data[604],
                             in_data[769]};
    
    wire lut_2167_out = lut_2167_table[lut_2167_select];
    
    generate
    if ( USE_REG ) begin : ff_2167
        reg   lut_2167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2167_ff <= lut_2167_out;
            end
        end
        
        assign out_data[2167] = lut_2167_ff;
    end
    else begin : no_ff_2167
        assign out_data[2167] = lut_2167_out;
    end
    endgenerate
    
    
    
    // LUT : 2168
    wire [63:0] lut_2168_table = 64'b0011001100110011000000000000000000000000001100110000000000000000;
    wire [5:0] lut_2168_select = {
                             in_data[185],
                             in_data[181],
                             in_data[161],
                             in_data[667],
                             in_data[683],
                             in_data[731]};
    
    wire lut_2168_out = lut_2168_table[lut_2168_select];
    
    generate
    if ( USE_REG ) begin : ff_2168
        reg   lut_2168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2168_ff <= lut_2168_out;
            end
        end
        
        assign out_data[2168] = lut_2168_ff;
    end
    else begin : no_ff_2168
        assign out_data[2168] = lut_2168_out;
    end
    endgenerate
    
    
    
    // LUT : 2169
    wire [63:0] lut_2169_table = 64'b0000000000000000100000001100000000001111000011110000111100001111;
    wire [5:0] lut_2169_select = {
                             in_data[359],
                             in_data[617],
                             in_data[280],
                             in_data[273],
                             in_data[722],
                             in_data[755]};
    
    wire lut_2169_out = lut_2169_table[lut_2169_select];
    
    generate
    if ( USE_REG ) begin : ff_2169
        reg   lut_2169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2169_ff <= lut_2169_out;
            end
        end
        
        assign out_data[2169] = lut_2169_ff;
    end
    else begin : no_ff_2169
        assign out_data[2169] = lut_2169_out;
    end
    endgenerate
    
    
    
    // LUT : 2170
    wire [63:0] lut_2170_table = 64'b1111111110001000111111111100110011111111110011001111111111001100;
    wire [5:0] lut_2170_select = {
                             in_data[725],
                             in_data[733],
                             in_data[678],
                             in_data[758],
                             in_data[318],
                             in_data[589]};
    
    wire lut_2170_out = lut_2170_table[lut_2170_select];
    
    generate
    if ( USE_REG ) begin : ff_2170
        reg   lut_2170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2170_ff <= lut_2170_out;
            end
        end
        
        assign out_data[2170] = lut_2170_ff;
    end
    else begin : no_ff_2170
        assign out_data[2170] = lut_2170_out;
    end
    endgenerate
    
    
    
    // LUT : 2171
    wire [63:0] lut_2171_table = 64'b0000010100000000000000000000000000001111000011110000111100001111;
    wire [5:0] lut_2171_select = {
                             in_data[119],
                             in_data[244],
                             in_data[79],
                             in_data[595],
                             in_data[585],
                             in_data[21]};
    
    wire lut_2171_out = lut_2171_table[lut_2171_select];
    
    generate
    if ( USE_REG ) begin : ff_2171
        reg   lut_2171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2171_ff <= lut_2171_out;
            end
        end
        
        assign out_data[2171] = lut_2171_ff;
    end
    else begin : no_ff_2171
        assign out_data[2171] = lut_2171_out;
    end
    endgenerate
    
    
    
    // LUT : 2172
    wire [63:0] lut_2172_table = 64'b0011001100110011001100110011001101110011001100110111001100110011;
    wire [5:0] lut_2172_select = {
                             in_data[613],
                             in_data[18],
                             in_data[677],
                             in_data[746],
                             in_data[547],
                             in_data[524]};
    
    wire lut_2172_out = lut_2172_table[lut_2172_select];
    
    generate
    if ( USE_REG ) begin : ff_2172
        reg   lut_2172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2172_ff <= lut_2172_out;
            end
        end
        
        assign out_data[2172] = lut_2172_ff;
    end
    else begin : no_ff_2172
        assign out_data[2172] = lut_2172_out;
    end
    endgenerate
    
    
    
    // LUT : 2173
    wire [63:0] lut_2173_table = 64'b0000000000000000101011111110111100000000000000001111111111101111;
    wire [5:0] lut_2173_select = {
                             in_data[391],
                             in_data[567],
                             in_data[448],
                             in_data[272],
                             in_data[698],
                             in_data[686]};
    
    wire lut_2173_out = lut_2173_table[lut_2173_select];
    
    generate
    if ( USE_REG ) begin : ff_2173
        reg   lut_2173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2173_ff <= lut_2173_out;
            end
        end
        
        assign out_data[2173] = lut_2173_ff;
    end
    else begin : no_ff_2173
        assign out_data[2173] = lut_2173_out;
    end
    endgenerate
    
    
    
    // LUT : 2174
    wire [63:0] lut_2174_table = 64'b0000000010001111000000000000000010001111111111110000000000001110;
    wire [5:0] lut_2174_select = {
                             in_data[397],
                             in_data[682],
                             in_data[362],
                             in_data[768],
                             in_data[675],
                             in_data[107]};
    
    wire lut_2174_out = lut_2174_table[lut_2174_select];
    
    generate
    if ( USE_REG ) begin : ff_2174
        reg   lut_2174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2174_ff <= lut_2174_out;
            end
        end
        
        assign out_data[2174] = lut_2174_ff;
    end
    else begin : no_ff_2174
        assign out_data[2174] = lut_2174_out;
    end
    endgenerate
    
    
    
    // LUT : 2175
    wire [63:0] lut_2175_table = 64'b0000000000000000001100000010000000000000000000001011001000110010;
    wire [5:0] lut_2175_select = {
                             in_data[367],
                             in_data[583],
                             in_data[8],
                             in_data[513],
                             in_data[739],
                             in_data[66]};
    
    wire lut_2175_out = lut_2175_table[lut_2175_select];
    
    generate
    if ( USE_REG ) begin : ff_2175
        reg   lut_2175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2175_ff <= lut_2175_out;
            end
        end
        
        assign out_data[2175] = lut_2175_ff;
    end
    else begin : no_ff_2175
        assign out_data[2175] = lut_2175_out;
    end
    endgenerate
    
    
    
    // LUT : 2176
    wire [63:0] lut_2176_table = 64'b1111001011110010111100101111001011111111111111111111001111110011;
    wire [5:0] lut_2176_select = {
                             in_data[151],
                             in_data[212],
                             in_data[46],
                             in_data[164],
                             in_data[573],
                             in_data[236]};
    
    wire lut_2176_out = lut_2176_table[lut_2176_select];
    
    generate
    if ( USE_REG ) begin : ff_2176
        reg   lut_2176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2176_ff <= lut_2176_out;
            end
        end
        
        assign out_data[2176] = lut_2176_ff;
    end
    else begin : no_ff_2176
        assign out_data[2176] = lut_2176_out;
    end
    endgenerate
    
    
    
    // LUT : 2177
    wire [63:0] lut_2177_table = 64'b0001001101110111000100010001000101110111011101010001000100010001;
    wire [5:0] lut_2177_select = {
                             in_data[554],
                             in_data[490],
                             in_data[40],
                             in_data[762],
                             in_data[400],
                             in_data[428]};
    
    wire lut_2177_out = lut_2177_table[lut_2177_select];
    
    generate
    if ( USE_REG ) begin : ff_2177
        reg   lut_2177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2177_ff <= lut_2177_out;
            end
        end
        
        assign out_data[2177] = lut_2177_ff;
    end
    else begin : no_ff_2177
        assign out_data[2177] = lut_2177_out;
    end
    endgenerate
    
    
    
    // LUT : 2178
    wire [63:0] lut_2178_table = 64'b1111111111001111111111111100111100000000110011000000000011001100;
    wire [5:0] lut_2178_select = {
                             in_data[261],
                             in_data[253],
                             in_data[369],
                             in_data[446],
                             in_data[342],
                             in_data[392]};
    
    wire lut_2178_out = lut_2178_table[lut_2178_select];
    
    generate
    if ( USE_REG ) begin : ff_2178
        reg   lut_2178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2178_ff <= lut_2178_out;
            end
        end
        
        assign out_data[2178] = lut_2178_ff;
    end
    else begin : no_ff_2178
        assign out_data[2178] = lut_2178_out;
    end
    endgenerate
    
    
    
    // LUT : 2179
    wire [63:0] lut_2179_table = 64'b0000000011000000000000000000000000001000110011000000100011001100;
    wire [5:0] lut_2179_select = {
                             in_data[690],
                             in_data[199],
                             in_data[153],
                             in_data[364],
                             in_data[601],
                             in_data[742]};
    
    wire lut_2179_out = lut_2179_table[lut_2179_select];
    
    generate
    if ( USE_REG ) begin : ff_2179
        reg   lut_2179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2179_ff <= lut_2179_out;
            end
        end
        
        assign out_data[2179] = lut_2179_ff;
    end
    else begin : no_ff_2179
        assign out_data[2179] = lut_2179_out;
    end
    endgenerate
    
    
    
    // LUT : 2180
    wire [63:0] lut_2180_table = 64'b1100110000000000111011110000000011111111000000001111111100000000;
    wire [5:0] lut_2180_select = {
                             in_data[534],
                             in_data[282],
                             in_data[370],
                             in_data[584],
                             in_data[91],
                             in_data[281]};
    
    wire lut_2180_out = lut_2180_table[lut_2180_select];
    
    generate
    if ( USE_REG ) begin : ff_2180
        reg   lut_2180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2180_ff <= lut_2180_out;
            end
        end
        
        assign out_data[2180] = lut_2180_ff;
    end
    else begin : no_ff_2180
        assign out_data[2180] = lut_2180_out;
    end
    endgenerate
    
    
    
    // LUT : 2181
    wire [63:0] lut_2181_table = 64'b1111111111111111111111111111000011111111111111111111111111110000;
    wire [5:0] lut_2181_select = {
                             in_data[284],
                             in_data[719],
                             in_data[296],
                             in_data[340],
                             in_data[449],
                             in_data[109]};
    
    wire lut_2181_out = lut_2181_table[lut_2181_select];
    
    generate
    if ( USE_REG ) begin : ff_2181
        reg   lut_2181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2181_ff <= lut_2181_out;
            end
        end
        
        assign out_data[2181] = lut_2181_ff;
    end
    else begin : no_ff_2181
        assign out_data[2181] = lut_2181_out;
    end
    endgenerate
    
    
    
    // LUT : 2182
    wire [63:0] lut_2182_table = 64'b0000010100000101000001010000010100000001000000010000010100000001;
    wire [5:0] lut_2182_select = {
                             in_data[42],
                             in_data[25],
                             in_data[444],
                             in_data[527],
                             in_data[108],
                             in_data[162]};
    
    wire lut_2182_out = lut_2182_table[lut_2182_select];
    
    generate
    if ( USE_REG ) begin : ff_2182
        reg   lut_2182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2182_ff <= lut_2182_out;
            end
        end
        
        assign out_data[2182] = lut_2182_ff;
    end
    else begin : no_ff_2182
        assign out_data[2182] = lut_2182_out;
    end
    endgenerate
    
    
    
    // LUT : 2183
    wire [63:0] lut_2183_table = 64'b0000000000000000000011110000000000001111000011110000111100001111;
    wire [5:0] lut_2183_select = {
                             in_data[489],
                             in_data[395],
                             in_data[502],
                             in_data[629],
                             in_data[533],
                             in_data[753]};
    
    wire lut_2183_out = lut_2183_table[lut_2183_select];
    
    generate
    if ( USE_REG ) begin : ff_2183
        reg   lut_2183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2183_ff <= lut_2183_out;
            end
        end
        
        assign out_data[2183] = lut_2183_ff;
    end
    else begin : no_ff_2183
        assign out_data[2183] = lut_2183_out;
    end
    endgenerate
    
    
    
    // LUT : 2184
    wire [63:0] lut_2184_table = 64'b0000111100001111000011110000111100001111000011110000111100001101;
    wire [5:0] lut_2184_select = {
                             in_data[776],
                             in_data[712],
                             in_data[777],
                             in_data[264],
                             in_data[780],
                             in_data[233]};
    
    wire lut_2184_out = lut_2184_table[lut_2184_select];
    
    generate
    if ( USE_REG ) begin : ff_2184
        reg   lut_2184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2184_ff <= lut_2184_out;
            end
        end
        
        assign out_data[2184] = lut_2184_ff;
    end
    else begin : no_ff_2184
        assign out_data[2184] = lut_2184_out;
    end
    endgenerate
    
    
    
    // LUT : 2185
    wire [63:0] lut_2185_table = 64'b1101110111111111000000001100110000000000010001000000000011011100;
    wire [5:0] lut_2185_select = {
                             in_data[346],
                             in_data[433],
                             in_data[649],
                             in_data[748],
                             in_data[221],
                             in_data[611]};
    
    wire lut_2185_out = lut_2185_table[lut_2185_select];
    
    generate
    if ( USE_REG ) begin : ff_2185
        reg   lut_2185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2185_ff <= lut_2185_out;
            end
        end
        
        assign out_data[2185] = lut_2185_ff;
    end
    else begin : no_ff_2185
        assign out_data[2185] = lut_2185_out;
    end
    endgenerate
    
    
    
    // LUT : 2186
    wire [63:0] lut_2186_table = 64'b1100111100000000100011110000000011111111000000001110111100000000;
    wire [5:0] lut_2186_select = {
                             in_data[130],
                             in_data[723],
                             in_data[382],
                             in_data[664],
                             in_data[424],
                             in_data[749]};
    
    wire lut_2186_out = lut_2186_table[lut_2186_select];
    
    generate
    if ( USE_REG ) begin : ff_2186
        reg   lut_2186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2186_ff <= lut_2186_out;
            end
        end
        
        assign out_data[2186] = lut_2186_ff;
    end
    else begin : no_ff_2186
        assign out_data[2186] = lut_2186_out;
    end
    endgenerate
    
    
    
    // LUT : 2187
    wire [63:0] lut_2187_table = 64'b0000111100001110000011110000111111111010111100101111101011110000;
    wire [5:0] lut_2187_select = {
                             in_data[320],
                             in_data[7],
                             in_data[50],
                             in_data[315],
                             in_data[219],
                             in_data[80]};
    
    wire lut_2187_out = lut_2187_table[lut_2187_select];
    
    generate
    if ( USE_REG ) begin : ff_2187
        reg   lut_2187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2187_ff <= lut_2187_out;
            end
        end
        
        assign out_data[2187] = lut_2187_ff;
    end
    else begin : no_ff_2187
        assign out_data[2187] = lut_2187_out;
    end
    endgenerate
    
    
    
    // LUT : 2188
    wire [63:0] lut_2188_table = 64'b1111000011111010111111111111101011110000101010101111101010101010;
    wire [5:0] lut_2188_select = {
                             in_data[535],
                             in_data[415],
                             in_data[457],
                             in_data[407],
                             in_data[557],
                             in_data[406]};
    
    wire lut_2188_out = lut_2188_table[lut_2188_select];
    
    generate
    if ( USE_REG ) begin : ff_2188
        reg   lut_2188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2188_ff <= lut_2188_out;
            end
        end
        
        assign out_data[2188] = lut_2188_ff;
    end
    else begin : no_ff_2188
        assign out_data[2188] = lut_2188_out;
    end
    endgenerate
    
    
    
    // LUT : 2189
    wire [63:0] lut_2189_table = 64'b0000000000000100011100011111000000000100100001000111000111110100;
    wire [5:0] lut_2189_select = {
                             in_data[39],
                             in_data[431],
                             in_data[207],
                             in_data[351],
                             in_data[345],
                             in_data[471]};
    
    wire lut_2189_out = lut_2189_table[lut_2189_select];
    
    generate
    if ( USE_REG ) begin : ff_2189
        reg   lut_2189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2189_ff <= lut_2189_out;
            end
        end
        
        assign out_data[2189] = lut_2189_ff;
    end
    else begin : no_ff_2189
        assign out_data[2189] = lut_2189_out;
    end
    endgenerate
    
    
    
    // LUT : 2190
    wire [63:0] lut_2190_table = 64'b0010101011111111101010101111111100000000111111110000000011101110;
    wire [5:0] lut_2190_select = {
                             in_data[217],
                             in_data[378],
                             in_data[210],
                             in_data[559],
                             in_data[636],
                             in_data[491]};
    
    wire lut_2190_out = lut_2190_table[lut_2190_select];
    
    generate
    if ( USE_REG ) begin : ff_2190
        reg   lut_2190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2190_ff <= lut_2190_out;
            end
        end
        
        assign out_data[2190] = lut_2190_ff;
    end
    else begin : no_ff_2190
        assign out_data[2190] = lut_2190_out;
    end
    endgenerate
    
    
    
    // LUT : 2191
    wire [63:0] lut_2191_table = 64'b1110111010101010111011101010101011101110101010101110111010101010;
    wire [5:0] lut_2191_select = {
                             in_data[530],
                             in_data[363],
                             in_data[631],
                             in_data[143],
                             in_data[497],
                             in_data[269]};
    
    wire lut_2191_out = lut_2191_table[lut_2191_select];
    
    generate
    if ( USE_REG ) begin : ff_2191
        reg   lut_2191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2191_ff <= lut_2191_out;
            end
        end
        
        assign out_data[2191] = lut_2191_ff;
    end
    else begin : no_ff_2191
        assign out_data[2191] = lut_2191_out;
    end
    endgenerate
    
    
    
    // LUT : 2192
    wire [63:0] lut_2192_table = 64'b1010101010111011101010101011101110101010101010101010101010101010;
    wire [5:0] lut_2192_select = {
                             in_data[721],
                             in_data[2],
                             in_data[188],
                             in_data[67],
                             in_data[705],
                             in_data[398]};
    
    wire lut_2192_out = lut_2192_table[lut_2192_select];
    
    generate
    if ( USE_REG ) begin : ff_2192
        reg   lut_2192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2192_ff <= lut_2192_out;
            end
        end
        
        assign out_data[2192] = lut_2192_ff;
    end
    else begin : no_ff_2192
        assign out_data[2192] = lut_2192_out;
    end
    endgenerate
    
    
    
    // LUT : 2193
    wire [63:0] lut_2193_table = 64'b0010001011111111000000001111111100100010111111110000000000001110;
    wire [5:0] lut_2193_select = {
                             in_data[577],
                             in_data[328],
                             in_data[403],
                             in_data[562],
                             in_data[688],
                             in_data[292]};
    
    wire lut_2193_out = lut_2193_table[lut_2193_select];
    
    generate
    if ( USE_REG ) begin : ff_2193
        reg   lut_2193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2193_ff <= lut_2193_out;
            end
        end
        
        assign out_data[2193] = lut_2193_ff;
    end
    else begin : no_ff_2193
        assign out_data[2193] = lut_2193_out;
    end
    endgenerate
    
    
    
    // LUT : 2194
    wire [63:0] lut_2194_table = 64'b1110111100000100111011111000111111101111000001011110111110001111;
    wire [5:0] lut_2194_select = {
                             in_data[476],
                             in_data[322],
                             in_data[555],
                             in_data[247],
                             in_data[528],
                             in_data[243]};
    
    wire lut_2194_out = lut_2194_table[lut_2194_select];
    
    generate
    if ( USE_REG ) begin : ff_2194
        reg   lut_2194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2194_ff <= lut_2194_out;
            end
        end
        
        assign out_data[2194] = lut_2194_ff;
    end
    else begin : no_ff_2194
        assign out_data[2194] = lut_2194_out;
    end
    endgenerate
    
    
    
    // LUT : 2195
    wire [63:0] lut_2195_table = 64'b1111110111111111000100010001000110111001111111110001000000010001;
    wire [5:0] lut_2195_select = {
                             in_data[53],
                             in_data[434],
                             in_data[355],
                             in_data[669],
                             in_data[241],
                             in_data[288]};
    
    wire lut_2195_out = lut_2195_table[lut_2195_select];
    
    generate
    if ( USE_REG ) begin : ff_2195
        reg   lut_2195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2195_ff <= lut_2195_out;
            end
        end
        
        assign out_data[2195] = lut_2195_ff;
    end
    else begin : no_ff_2195
        assign out_data[2195] = lut_2195_out;
    end
    endgenerate
    
    
    
    // LUT : 2196
    wire [63:0] lut_2196_table = 64'b1111111111111111000000000000010011111111111111111111111111111111;
    wire [5:0] lut_2196_select = {
                             in_data[437],
                             in_data[255],
                             in_data[87],
                             in_data[168],
                             in_data[154],
                             in_data[699]};
    
    wire lut_2196_out = lut_2196_table[lut_2196_select];
    
    generate
    if ( USE_REG ) begin : ff_2196
        reg   lut_2196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2196_ff <= lut_2196_out;
            end
        end
        
        assign out_data[2196] = lut_2196_ff;
    end
    else begin : no_ff_2196
        assign out_data[2196] = lut_2196_out;
    end
    endgenerate
    
    
    
    // LUT : 2197
    wire [63:0] lut_2197_table = 64'b0000000011001100111111111100111110111111001111110011001100000000;
    wire [5:0] lut_2197_select = {
                             in_data[543],
                             in_data[483],
                             in_data[283],
                             in_data[6],
                             in_data[182],
                             in_data[727]};
    
    wire lut_2197_out = lut_2197_table[lut_2197_select];
    
    generate
    if ( USE_REG ) begin : ff_2197
        reg   lut_2197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2197_ff <= lut_2197_out;
            end
        end
        
        assign out_data[2197] = lut_2197_ff;
    end
    else begin : no_ff_2197
        assign out_data[2197] = lut_2197_out;
    end
    endgenerate
    
    
    
    // LUT : 2198
    wire [63:0] lut_2198_table = 64'b0000000011111111111111111111111100000000000000000000000011111111;
    wire [5:0] lut_2198_select = {
                             in_data[472],
                             in_data[285],
                             in_data[356],
                             in_data[532],
                             in_data[334],
                             in_data[778]};
    
    wire lut_2198_out = lut_2198_table[lut_2198_select];
    
    generate
    if ( USE_REG ) begin : ff_2198
        reg   lut_2198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2198_ff <= lut_2198_out;
            end
        end
        
        assign out_data[2198] = lut_2198_ff;
    end
    else begin : no_ff_2198
        assign out_data[2198] = lut_2198_out;
    end
    endgenerate
    
    
    
    // LUT : 2199
    wire [63:0] lut_2199_table = 64'b0000000000000000111111111111111100000000000000001110111111111111;
    wire [5:0] lut_2199_select = {
                             in_data[250],
                             in_data[150],
                             in_data[15],
                             in_data[413],
                             in_data[339],
                             in_data[306]};
    
    wire lut_2199_out = lut_2199_table[lut_2199_select];
    
    generate
    if ( USE_REG ) begin : ff_2199
        reg   lut_2199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2199_ff <= lut_2199_out;
            end
        end
        
        assign out_data[2199] = lut_2199_ff;
    end
    else begin : no_ff_2199
        assign out_data[2199] = lut_2199_out;
    end
    endgenerate
    
    
    
    // LUT : 2200
    wire [63:0] lut_2200_table = 64'b1011000010111010001100001011101010110000101110100011000010111010;
    wire [5:0] lut_2200_select = {
                             in_data[366],
                             in_data[475],
                             in_data[330],
                             in_data[602],
                             in_data[135],
                             in_data[177]};
    
    wire lut_2200_out = lut_2200_table[lut_2200_select];
    
    generate
    if ( USE_REG ) begin : ff_2200
        reg   lut_2200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2200_ff <= lut_2200_out;
            end
        end
        
        assign out_data[2200] = lut_2200_ff;
    end
    else begin : no_ff_2200
        assign out_data[2200] = lut_2200_out;
    end
    endgenerate
    
    
    
    // LUT : 2201
    wire [63:0] lut_2201_table = 64'b0000000101010101000000010101010100000101000001010000010100000001;
    wire [5:0] lut_2201_select = {
                             in_data[576],
                             in_data[4],
                             in_data[581],
                             in_data[599],
                             in_data[170],
                             in_data[123]};
    
    wire lut_2201_out = lut_2201_table[lut_2201_select];
    
    generate
    if ( USE_REG ) begin : ff_2201
        reg   lut_2201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2201_ff <= lut_2201_out;
            end
        end
        
        assign out_data[2201] = lut_2201_ff;
    end
    else begin : no_ff_2201
        assign out_data[2201] = lut_2201_out;
    end
    endgenerate
    
    
    
    // LUT : 2202
    wire [63:0] lut_2202_table = 64'b1111111111111111111111111111111101010100010101001101010011010100;
    wire [5:0] lut_2202_select = {
                             in_data[624],
                             in_data[672],
                             in_data[136],
                             in_data[347],
                             in_data[312],
                             in_data[101]};
    
    wire lut_2202_out = lut_2202_table[lut_2202_select];
    
    generate
    if ( USE_REG ) begin : ff_2202
        reg   lut_2202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2202_ff <= lut_2202_out;
            end
        end
        
        assign out_data[2202] = lut_2202_ff;
    end
    else begin : no_ff_2202
        assign out_data[2202] = lut_2202_out;
    end
    endgenerate
    
    
    
    // LUT : 2203
    wire [63:0] lut_2203_table = 64'b0000010000001100000000000000000011001101110011110000110000001100;
    wire [5:0] lut_2203_select = {
                             in_data[404],
                             in_data[71],
                             in_data[474],
                             in_data[650],
                             in_data[263],
                             in_data[642]};
    
    wire lut_2203_out = lut_2203_table[lut_2203_select];
    
    generate
    if ( USE_REG ) begin : ff_2203
        reg   lut_2203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2203_ff <= lut_2203_out;
            end
        end
        
        assign out_data[2203] = lut_2203_ff;
    end
    else begin : no_ff_2203
        assign out_data[2203] = lut_2203_out;
    end
    endgenerate
    
    
    
    // LUT : 2204
    wire [63:0] lut_2204_table = 64'b0010001100100011000000000000000011111111111011101100110011001100;
    wire [5:0] lut_2204_select = {
                             in_data[662],
                             in_data[520],
                             in_data[117],
                             in_data[13],
                             in_data[516],
                             in_data[390]};
    
    wire lut_2204_out = lut_2204_table[lut_2204_select];
    
    generate
    if ( USE_REG ) begin : ff_2204
        reg   lut_2204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2204_ff <= lut_2204_out;
            end
        end
        
        assign out_data[2204] = lut_2204_ff;
    end
    else begin : no_ff_2204
        assign out_data[2204] = lut_2204_out;
    end
    endgenerate
    
    
    
    // LUT : 2205
    wire [63:0] lut_2205_table = 64'b1111111111111111101011110000101111111111111111111010111100001111;
    wire [5:0] lut_2205_select = {
                             in_data[591],
                             in_data[498],
                             in_data[445],
                             in_data[515],
                             in_data[618],
                             in_data[72]};
    
    wire lut_2205_out = lut_2205_table[lut_2205_select];
    
    generate
    if ( USE_REG ) begin : ff_2205
        reg   lut_2205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2205_ff <= lut_2205_out;
            end
        end
        
        assign out_data[2205] = lut_2205_ff;
    end
    else begin : no_ff_2205
        assign out_data[2205] = lut_2205_out;
    end
    endgenerate
    
    
    
    // LUT : 2206
    wire [63:0] lut_2206_table = 64'b1111111111110000111111111111000011111100111100001111111111110000;
    wire [5:0] lut_2206_select = {
                             in_data[60],
                             in_data[365],
                             in_data[603],
                             in_data[432],
                             in_data[561],
                             in_data[30]};
    
    wire lut_2206_out = lut_2206_table[lut_2206_select];
    
    generate
    if ( USE_REG ) begin : ff_2206
        reg   lut_2206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2206_ff <= lut_2206_out;
            end
        end
        
        assign out_data[2206] = lut_2206_ff;
    end
    else begin : no_ff_2206
        assign out_data[2206] = lut_2206_out;
    end
    endgenerate
    
    
    
    // LUT : 2207
    wire [63:0] lut_2207_table = 64'b1111110011011100111111001101110111111000110111011111110011011101;
    wire [5:0] lut_2207_select = {
                             in_data[222],
                             in_data[36],
                             in_data[487],
                             in_data[417],
                             in_data[454],
                             in_data[146]};
    
    wire lut_2207_out = lut_2207_table[lut_2207_select];
    
    generate
    if ( USE_REG ) begin : ff_2207
        reg   lut_2207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2207_ff <= lut_2207_out;
            end
        end
        
        assign out_data[2207] = lut_2207_ff;
    end
    else begin : no_ff_2207
        assign out_data[2207] = lut_2207_out;
    end
    endgenerate
    
    
    
    // LUT : 2208
    wire [63:0] lut_2208_table = 64'b1100111111001100000000110000110011001111110011000000001100001100;
    wire [5:0] lut_2208_select = {
                             in_data[616],
                             in_data[623],
                             in_data[605],
                             in_data[248],
                             in_data[552],
                             in_data[141]};
    
    wire lut_2208_out = lut_2208_table[lut_2208_select];
    
    generate
    if ( USE_REG ) begin : ff_2208
        reg   lut_2208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2208_ff <= lut_2208_out;
            end
        end
        
        assign out_data[2208] = lut_2208_ff;
    end
    else begin : no_ff_2208
        assign out_data[2208] = lut_2208_out;
    end
    endgenerate
    
    
    
    // LUT : 2209
    wire [63:0] lut_2209_table = 64'b0000000000000000000000000000001100000000000000000000000000000011;
    wire [5:0] lut_2209_select = {
                             in_data[259],
                             in_data[509],
                             in_data[313],
                             in_data[387],
                             in_data[173],
                             in_data[172]};
    
    wire lut_2209_out = lut_2209_table[lut_2209_select];
    
    generate
    if ( USE_REG ) begin : ff_2209
        reg   lut_2209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2209_ff <= lut_2209_out;
            end
        end
        
        assign out_data[2209] = lut_2209_ff;
    end
    else begin : no_ff_2209
        assign out_data[2209] = lut_2209_out;
    end
    endgenerate
    
    
    
    // LUT : 2210
    wire [63:0] lut_2210_table = 64'b0000000100000000111111111101111100000011000000001111111111111111;
    wire [5:0] lut_2210_select = {
                             in_data[721],
                             in_data[435],
                             in_data[633],
                             in_data[131],
                             in_data[401],
                             in_data[24]};
    
    wire lut_2210_out = lut_2210_table[lut_2210_select];
    
    generate
    if ( USE_REG ) begin : ff_2210
        reg   lut_2210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2210_ff <= lut_2210_out;
            end
        end
        
        assign out_data[2210] = lut_2210_ff;
    end
    else begin : no_ff_2210
        assign out_data[2210] = lut_2210_out;
    end
    endgenerate
    
    
    
    // LUT : 2211
    wire [63:0] lut_2211_table = 64'b1010101010101111000010000000101010101010111111111111000011111010;
    wire [5:0] lut_2211_select = {
                             in_data[635],
                             in_data[190],
                             in_data[157],
                             in_data[323],
                             in_data[703],
                             in_data[192]};
    
    wire lut_2211_out = lut_2211_table[lut_2211_select];
    
    generate
    if ( USE_REG ) begin : ff_2211
        reg   lut_2211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2211_ff <= lut_2211_out;
            end
        end
        
        assign out_data[2211] = lut_2211_ff;
    end
    else begin : no_ff_2211
        assign out_data[2211] = lut_2211_out;
    end
    endgenerate
    
    
    
    // LUT : 2212
    wire [63:0] lut_2212_table = 64'b1110000011000000111000001111000011110000111111111111000011111111;
    wire [5:0] lut_2212_select = {
                             in_data[487],
                             in_data[79],
                             in_data[652],
                             in_data[342],
                             in_data[68],
                             in_data[731]};
    
    wire lut_2212_out = lut_2212_table[lut_2212_select];
    
    generate
    if ( USE_REG ) begin : ff_2212
        reg   lut_2212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2212_ff <= lut_2212_out;
            end
        end
        
        assign out_data[2212] = lut_2212_ff;
    end
    else begin : no_ff_2212
        assign out_data[2212] = lut_2212_out;
    end
    endgenerate
    
    
    
    // LUT : 2213
    wire [63:0] lut_2213_table = 64'b1111111111111111100011110000110111111111111011111000111100001111;
    wire [5:0] lut_2213_select = {
                             in_data[15],
                             in_data[481],
                             in_data[171],
                             in_data[233],
                             in_data[104],
                             in_data[217]};
    
    wire lut_2213_out = lut_2213_table[lut_2213_select];
    
    generate
    if ( USE_REG ) begin : ff_2213
        reg   lut_2213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2213_ff <= lut_2213_out;
            end
        end
        
        assign out_data[2213] = lut_2213_ff;
    end
    else begin : no_ff_2213
        assign out_data[2213] = lut_2213_out;
    end
    endgenerate
    
    
    
    // LUT : 2214
    wire [63:0] lut_2214_table = 64'b0011011111111111000000000011000000110011111111110000000000100000;
    wire [5:0] lut_2214_select = {
                             in_data[733],
                             in_data[243],
                             in_data[63],
                             in_data[456],
                             in_data[597],
                             in_data[448]};
    
    wire lut_2214_out = lut_2214_table[lut_2214_select];
    
    generate
    if ( USE_REG ) begin : ff_2214
        reg   lut_2214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2214_ff <= lut_2214_out;
            end
        end
        
        assign out_data[2214] = lut_2214_ff;
    end
    else begin : no_ff_2214
        assign out_data[2214] = lut_2214_out;
    end
    endgenerate
    
    
    
    // LUT : 2215
    wire [63:0] lut_2215_table = 64'b1111101000101010000010100000101011111111111110111111101010101010;
    wire [5:0] lut_2215_select = {
                             in_data[317],
                             in_data[565],
                             in_data[74],
                             in_data[489],
                             in_data[730],
                             in_data[270]};
    
    wire lut_2215_out = lut_2215_table[lut_2215_select];
    
    generate
    if ( USE_REG ) begin : ff_2215
        reg   lut_2215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2215_ff <= lut_2215_out;
            end
        end
        
        assign out_data[2215] = lut_2215_ff;
    end
    else begin : no_ff_2215
        assign out_data[2215] = lut_2215_out;
    end
    endgenerate
    
    
    
    // LUT : 2216
    wire [63:0] lut_2216_table = 64'b0100010001001100010001000100010001000100010011000100010001000100;
    wire [5:0] lut_2216_select = {
                             in_data[141],
                             in_data[383],
                             in_data[92],
                             in_data[255],
                             in_data[627],
                             in_data[444]};
    
    wire lut_2216_out = lut_2216_table[lut_2216_select];
    
    generate
    if ( USE_REG ) begin : ff_2216
        reg   lut_2216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2216_ff <= lut_2216_out;
            end
        end
        
        assign out_data[2216] = lut_2216_ff;
    end
    else begin : no_ff_2216
        assign out_data[2216] = lut_2216_out;
    end
    endgenerate
    
    
    
    // LUT : 2217
    wire [63:0] lut_2217_table = 64'b1010111110101111000000000000010110101111101011110000000000000101;
    wire [5:0] lut_2217_select = {
                             in_data[196],
                             in_data[207],
                             in_data[594],
                             in_data[655],
                             in_data[670],
                             in_data[341]};
    
    wire lut_2217_out = lut_2217_table[lut_2217_select];
    
    generate
    if ( USE_REG ) begin : ff_2217
        reg   lut_2217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2217_ff <= lut_2217_out;
            end
        end
        
        assign out_data[2217] = lut_2217_ff;
    end
    else begin : no_ff_2217
        assign out_data[2217] = lut_2217_out;
    end
    endgenerate
    
    
    
    // LUT : 2218
    wire [63:0] lut_2218_table = 64'b0000010100000101000000000000000001011111010111110000000000000000;
    wire [5:0] lut_2218_select = {
                             in_data[151],
                             in_data[488],
                             in_data[31],
                             in_data[125],
                             in_data[34],
                             in_data[611]};
    
    wire lut_2218_out = lut_2218_table[lut_2218_select];
    
    generate
    if ( USE_REG ) begin : ff_2218
        reg   lut_2218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2218_ff <= lut_2218_out;
            end
        end
        
        assign out_data[2218] = lut_2218_ff;
    end
    else begin : no_ff_2218
        assign out_data[2218] = lut_2218_out;
    end
    endgenerate
    
    
    
    // LUT : 2219
    wire [63:0] lut_2219_table = 64'b1111111111011101111111111111111111000100000000001111111111111111;
    wire [5:0] lut_2219_select = {
                             in_data[119],
                             in_data[689],
                             in_data[43],
                             in_data[726],
                             in_data[222],
                             in_data[509]};
    
    wire lut_2219_out = lut_2219_table[lut_2219_select];
    
    generate
    if ( USE_REG ) begin : ff_2219
        reg   lut_2219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2219_ff <= lut_2219_out;
            end
        end
        
        assign out_data[2219] = lut_2219_ff;
    end
    else begin : no_ff_2219
        assign out_data[2219] = lut_2219_out;
    end
    endgenerate
    
    
    
    // LUT : 2220
    wire [63:0] lut_2220_table = 64'b0000000011110000000000000011000000000000111100000000000000110000;
    wire [5:0] lut_2220_select = {
                             in_data[449],
                             in_data[267],
                             in_data[556],
                             in_data[380],
                             in_data[388],
                             in_data[700]};
    
    wire lut_2220_out = lut_2220_table[lut_2220_select];
    
    generate
    if ( USE_REG ) begin : ff_2220
        reg   lut_2220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2220_ff <= lut_2220_out;
            end
        end
        
        assign out_data[2220] = lut_2220_ff;
    end
    else begin : no_ff_2220
        assign out_data[2220] = lut_2220_out;
    end
    endgenerate
    
    
    
    // LUT : 2221
    wire [63:0] lut_2221_table = 64'b0000000001010101000000000101010110000000111111111000100011111101;
    wire [5:0] lut_2221_select = {
                             in_data[324],
                             in_data[748],
                             in_data[378],
                             in_data[504],
                             in_data[554],
                             in_data[538]};
    
    wire lut_2221_out = lut_2221_table[lut_2221_select];
    
    generate
    if ( USE_REG ) begin : ff_2221
        reg   lut_2221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2221_ff <= lut_2221_out;
            end
        end
        
        assign out_data[2221] = lut_2221_ff;
    end
    else begin : no_ff_2221
        assign out_data[2221] = lut_2221_out;
    end
    endgenerate
    
    
    
    // LUT : 2222
    wire [63:0] lut_2222_table = 64'b1111111111111111100011001000110011111111111111111010101010101010;
    wire [5:0] lut_2222_select = {
                             in_data[289],
                             in_data[101],
                             in_data[20],
                             in_data[459],
                             in_data[482],
                             in_data[578]};
    
    wire lut_2222_out = lut_2222_table[lut_2222_select];
    
    generate
    if ( USE_REG ) begin : ff_2222
        reg   lut_2222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2222_ff <= lut_2222_out;
            end
        end
        
        assign out_data[2222] = lut_2222_ff;
    end
    else begin : no_ff_2222
        assign out_data[2222] = lut_2222_out;
    end
    endgenerate
    
    
    
    // LUT : 2223
    wire [63:0] lut_2223_table = 64'b1111111111111111111111111111111111111111111011101111111111101110;
    wire [5:0] lut_2223_select = {
                             in_data[362],
                             in_data[617],
                             in_data[135],
                             in_data[771],
                             in_data[262],
                             in_data[163]};
    
    wire lut_2223_out = lut_2223_table[lut_2223_select];
    
    generate
    if ( USE_REG ) begin : ff_2223
        reg   lut_2223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2223_ff <= lut_2223_out;
            end
        end
        
        assign out_data[2223] = lut_2223_ff;
    end
    else begin : no_ff_2223
        assign out_data[2223] = lut_2223_out;
    end
    endgenerate
    
    
    
    // LUT : 2224
    wire [63:0] lut_2224_table = 64'b1000111010001111111111111110111110001110000011111111111110101111;
    wire [5:0] lut_2224_select = {
                             in_data[14],
                             in_data[600],
                             in_data[431],
                             in_data[269],
                             in_data[678],
                             in_data[332]};
    
    wire lut_2224_out = lut_2224_table[lut_2224_select];
    
    generate
    if ( USE_REG ) begin : ff_2224
        reg   lut_2224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2224_ff <= lut_2224_out;
            end
        end
        
        assign out_data[2224] = lut_2224_ff;
    end
    else begin : no_ff_2224
        assign out_data[2224] = lut_2224_out;
    end
    endgenerate
    
    
    
    // LUT : 2225
    wire [63:0] lut_2225_table = 64'b1111111111111111111111001111111111111100111111111100000011111111;
    wire [5:0] lut_2225_select = {
                             in_data[591],
                             in_data[127],
                             in_data[379],
                             in_data[256],
                             in_data[390],
                             in_data[145]};
    
    wire lut_2225_out = lut_2225_table[lut_2225_select];
    
    generate
    if ( USE_REG ) begin : ff_2225
        reg   lut_2225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2225_ff <= lut_2225_out;
            end
        end
        
        assign out_data[2225] = lut_2225_ff;
    end
    else begin : no_ff_2225
        assign out_data[2225] = lut_2225_out;
    end
    endgenerate
    
    
    
    // LUT : 2226
    wire [63:0] lut_2226_table = 64'b0001000101110111000000000000000001010001011101110000000000000000;
    wire [5:0] lut_2226_select = {
                             in_data[675],
                             in_data[549],
                             in_data[299],
                             in_data[767],
                             in_data[276],
                             in_data[311]};
    
    wire lut_2226_out = lut_2226_table[lut_2226_select];
    
    generate
    if ( USE_REG ) begin : ff_2226
        reg   lut_2226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2226_ff <= lut_2226_out;
            end
        end
        
        assign out_data[2226] = lut_2226_ff;
    end
    else begin : no_ff_2226
        assign out_data[2226] = lut_2226_out;
    end
    endgenerate
    
    
    
    // LUT : 2227
    wire [63:0] lut_2227_table = 64'b1111111111111110111111111111111011111111111100001111111111110000;
    wire [5:0] lut_2227_select = {
                             in_data[497],
                             in_data[9],
                             in_data[619],
                             in_data[156],
                             in_data[35],
                             in_data[697]};
    
    wire lut_2227_out = lut_2227_table[lut_2227_select];
    
    generate
    if ( USE_REG ) begin : ff_2227
        reg   lut_2227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2227_ff <= lut_2227_out;
            end
        end
        
        assign out_data[2227] = lut_2227_ff;
    end
    else begin : no_ff_2227
        assign out_data[2227] = lut_2227_out;
    end
    endgenerate
    
    
    
    // LUT : 2228
    wire [63:0] lut_2228_table = 64'b0011000100010001111100010001000110111011000000001011101100000000;
    wire [5:0] lut_2228_select = {
                             in_data[209],
                             in_data[503],
                             in_data[355],
                             in_data[186],
                             in_data[592],
                             in_data[657]};
    
    wire lut_2228_out = lut_2228_table[lut_2228_select];
    
    generate
    if ( USE_REG ) begin : ff_2228
        reg   lut_2228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2228_ff <= lut_2228_out;
            end
        end
        
        assign out_data[2228] = lut_2228_ff;
    end
    else begin : no_ff_2228
        assign out_data[2228] = lut_2228_out;
    end
    endgenerate
    
    
    
    // LUT : 2229
    wire [63:0] lut_2229_table = 64'b0000000000000000000011110000000000000000000000001111111111111111;
    wire [5:0] lut_2229_select = {
                             in_data[381],
                             in_data[414],
                             in_data[574],
                             in_data[226],
                             in_data[724],
                             in_data[62]};
    
    wire lut_2229_out = lut_2229_table[lut_2229_select];
    
    generate
    if ( USE_REG ) begin : ff_2229
        reg   lut_2229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2229_ff <= lut_2229_out;
            end
        end
        
        assign out_data[2229] = lut_2229_ff;
    end
    else begin : no_ff_2229
        assign out_data[2229] = lut_2229_out;
    end
    endgenerate
    
    
    
    // LUT : 2230
    wire [63:0] lut_2230_table = 64'b1100110011001100010001001100110011001100110011000100010011001100;
    wire [5:0] lut_2230_select = {
                             in_data[18],
                             in_data[551],
                             in_data[518],
                             in_data[589],
                             in_data[329],
                             in_data[708]};
    
    wire lut_2230_out = lut_2230_table[lut_2230_select];
    
    generate
    if ( USE_REG ) begin : ff_2230
        reg   lut_2230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2230_ff <= lut_2230_out;
            end
        end
        
        assign out_data[2230] = lut_2230_ff;
    end
    else begin : no_ff_2230
        assign out_data[2230] = lut_2230_out;
    end
    endgenerate
    
    
    
    // LUT : 2231
    wire [63:0] lut_2231_table = 64'b0101000011110101000000001111010100000000011101010000000001110101;
    wire [5:0] lut_2231_select = {
                             in_data[280],
                             in_data[98],
                             in_data[133],
                             in_data[593],
                             in_data[5],
                             in_data[387]};
    
    wire lut_2231_out = lut_2231_table[lut_2231_select];
    
    generate
    if ( USE_REG ) begin : ff_2231
        reg   lut_2231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2231_ff <= lut_2231_out;
            end
        end
        
        assign out_data[2231] = lut_2231_ff;
    end
    else begin : no_ff_2231
        assign out_data[2231] = lut_2231_out;
    end
    endgenerate
    
    
    
    // LUT : 2232
    wire [63:0] lut_2232_table = 64'b1110101011101110110010001100100011111111111011101100110011101110;
    wire [5:0] lut_2232_select = {
                             in_data[248],
                             in_data[344],
                             in_data[439],
                             in_data[279],
                             in_data[491],
                             in_data[536]};
    
    wire lut_2232_out = lut_2232_table[lut_2232_select];
    
    generate
    if ( USE_REG ) begin : ff_2232
        reg   lut_2232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2232_ff <= lut_2232_out;
            end
        end
        
        assign out_data[2232] = lut_2232_ff;
    end
    else begin : no_ff_2232
        assign out_data[2232] = lut_2232_out;
    end
    endgenerate
    
    
    
    // LUT : 2233
    wire [63:0] lut_2233_table = 64'b0100010001000100010001000100010001000100010001000100010001000100;
    wire [5:0] lut_2233_select = {
                             in_data[746],
                             in_data[662],
                             in_data[763],
                             in_data[28],
                             in_data[517],
                             in_data[330]};
    
    wire lut_2233_out = lut_2233_table[lut_2233_select];
    
    generate
    if ( USE_REG ) begin : ff_2233
        reg   lut_2233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2233_ff <= lut_2233_out;
            end
        end
        
        assign out_data[2233] = lut_2233_ff;
    end
    else begin : no_ff_2233
        assign out_data[2233] = lut_2233_out;
    end
    endgenerate
    
    
    
    // LUT : 2234
    wire [63:0] lut_2234_table = 64'b0000000000000000000000000000000011001100110011001100110011011100;
    wire [5:0] lut_2234_select = {
                             in_data[183],
                             in_data[224],
                             in_data[775],
                             in_data[272],
                             in_data[318],
                             in_data[142]};
    
    wire lut_2234_out = lut_2234_table[lut_2234_select];
    
    generate
    if ( USE_REG ) begin : ff_2234
        reg   lut_2234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2234_ff <= lut_2234_out;
            end
        end
        
        assign out_data[2234] = lut_2234_ff;
    end
    else begin : no_ff_2234
        assign out_data[2234] = lut_2234_out;
    end
    endgenerate
    
    
    
    // LUT : 2235
    wire [63:0] lut_2235_table = 64'b1111111111111111111111111111111111111111111110101111111111111010;
    wire [5:0] lut_2235_select = {
                             in_data[744],
                             in_data[359],
                             in_data[221],
                             in_data[707],
                             in_data[364],
                             in_data[628]};
    
    wire lut_2235_out = lut_2235_table[lut_2235_select];
    
    generate
    if ( USE_REG ) begin : ff_2235
        reg   lut_2235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2235_ff <= lut_2235_out;
            end
        end
        
        assign out_data[2235] = lut_2235_ff;
    end
    else begin : no_ff_2235
        assign out_data[2235] = lut_2235_out;
    end
    endgenerate
    
    
    
    // LUT : 2236
    wire [63:0] lut_2236_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_2236_select = {
                             in_data[258],
                             in_data[360],
                             in_data[144],
                             in_data[89],
                             in_data[615],
                             in_data[507]};
    
    wire lut_2236_out = lut_2236_table[lut_2236_select];
    
    generate
    if ( USE_REG ) begin : ff_2236
        reg   lut_2236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2236_ff <= lut_2236_out;
            end
        end
        
        assign out_data[2236] = lut_2236_ff;
    end
    else begin : no_ff_2236
        assign out_data[2236] = lut_2236_out;
    end
    endgenerate
    
    
    
    // LUT : 2237
    wire [63:0] lut_2237_table = 64'b1111110011111110111111111111111111110000111110001111110011111100;
    wire [5:0] lut_2237_select = {
                             in_data[120],
                             in_data[165],
                             in_data[282],
                             in_data[174],
                             in_data[423],
                             in_data[643]};
    
    wire lut_2237_out = lut_2237_table[lut_2237_select];
    
    generate
    if ( USE_REG ) begin : ff_2237
        reg   lut_2237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2237_ff <= lut_2237_out;
            end
        end
        
        assign out_data[2237] = lut_2237_ff;
    end
    else begin : no_ff_2237
        assign out_data[2237] = lut_2237_out;
    end
    endgenerate
    
    
    
    // LUT : 2238
    wire [63:0] lut_2238_table = 64'b1111111001000100111111111100110001000100010101010101110101010101;
    wire [5:0] lut_2238_select = {
                             in_data[440],
                             in_data[566],
                             in_data[580],
                             in_data[339],
                             in_data[219],
                             in_data[469]};
    
    wire lut_2238_out = lut_2238_table[lut_2238_select];
    
    generate
    if ( USE_REG ) begin : ff_2238
        reg   lut_2238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2238_ff <= lut_2238_out;
            end
        end
        
        assign out_data[2238] = lut_2238_ff;
    end
    else begin : no_ff_2238
        assign out_data[2238] = lut_2238_out;
    end
    endgenerate
    
    
    
    // LUT : 2239
    wire [63:0] lut_2239_table = 64'b1010111110101111000011110000111100111111101111110000101100001011;
    wire [5:0] lut_2239_select = {
                             in_data[19],
                             in_data[676],
                             in_data[738],
                             in_data[749],
                             in_data[585],
                             in_data[642]};
    
    wire lut_2239_out = lut_2239_table[lut_2239_select];
    
    generate
    if ( USE_REG ) begin : ff_2239
        reg   lut_2239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2239_ff <= lut_2239_out;
            end
        end
        
        assign out_data[2239] = lut_2239_ff;
    end
    else begin : no_ff_2239
        assign out_data[2239] = lut_2239_out;
    end
    endgenerate
    
    
    
    // LUT : 2240
    wire [63:0] lut_2240_table = 64'b0000101000001010010101010101010100001010000000100100010101010101;
    wire [5:0] lut_2240_select = {
                             in_data[776],
                             in_data[512],
                             in_data[666],
                             in_data[546],
                             in_data[69],
                             in_data[541]};
    
    wire lut_2240_out = lut_2240_table[lut_2240_select];
    
    generate
    if ( USE_REG ) begin : ff_2240
        reg   lut_2240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2240_ff <= lut_2240_out;
            end
        end
        
        assign out_data[2240] = lut_2240_ff;
    end
    else begin : no_ff_2240
        assign out_data[2240] = lut_2240_out;
    end
    endgenerate
    
    
    
    // LUT : 2241
    wire [63:0] lut_2241_table = 64'b1110110011101100111111101111111011101100111011001111111011101100;
    wire [5:0] lut_2241_select = {
                             in_data[117],
                             in_data[712],
                             in_data[65],
                             in_data[278],
                             in_data[493],
                             in_data[99]};
    
    wire lut_2241_out = lut_2241_table[lut_2241_select];
    
    generate
    if ( USE_REG ) begin : ff_2241
        reg   lut_2241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2241_ff <= lut_2241_out;
            end
        end
        
        assign out_data[2241] = lut_2241_ff;
    end
    else begin : no_ff_2241
        assign out_data[2241] = lut_2241_out;
    end
    endgenerate
    
    
    
    // LUT : 2242
    wire [63:0] lut_2242_table = 64'b1111111111111111111111111011111111111111111111111011101100110011;
    wire [5:0] lut_2242_select = {
                             in_data[528],
                             in_data[457],
                             in_data[223],
                             in_data[16],
                             in_data[434],
                             in_data[684]};
    
    wire lut_2242_out = lut_2242_table[lut_2242_select];
    
    generate
    if ( USE_REG ) begin : ff_2242
        reg   lut_2242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2242_ff <= lut_2242_out;
            end
        end
        
        assign out_data[2242] = lut_2242_ff;
    end
    else begin : no_ff_2242
        assign out_data[2242] = lut_2242_out;
    end
    endgenerate
    
    
    
    // LUT : 2243
    wire [63:0] lut_2243_table = 64'b0101000000001111010100000000111101010000000111110101000000001010;
    wire [5:0] lut_2243_select = {
                             in_data[44],
                             in_data[639],
                             in_data[564],
                             in_data[460],
                             in_data[252],
                             in_data[384]};
    
    wire lut_2243_out = lut_2243_table[lut_2243_select];
    
    generate
    if ( USE_REG ) begin : ff_2243
        reg   lut_2243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2243_ff <= lut_2243_out;
            end
        end
        
        assign out_data[2243] = lut_2243_ff;
    end
    else begin : no_ff_2243
        assign out_data[2243] = lut_2243_out;
    end
    endgenerate
    
    
    
    // LUT : 2244
    wire [63:0] lut_2244_table = 64'b1111010011110000111111111111001101010000011100001111111111110001;
    wire [5:0] lut_2244_select = {
                             in_data[772],
                             in_data[77],
                             in_data[468],
                             in_data[176],
                             in_data[350],
                             in_data[191]};
    
    wire lut_2244_out = lut_2244_table[lut_2244_select];
    
    generate
    if ( USE_REG ) begin : ff_2244
        reg   lut_2244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2244_ff <= lut_2244_out;
            end
        end
        
        assign out_data[2244] = lut_2244_ff;
    end
    else begin : no_ff_2244
        assign out_data[2244] = lut_2244_out;
    end
    endgenerate
    
    
    
    // LUT : 2245
    wire [63:0] lut_2245_table = 64'b1011001011111111101100101111111110100000101100111010000010110011;
    wire [5:0] lut_2245_select = {
                             in_data[331],
                             in_data[32],
                             in_data[305],
                             in_data[261],
                             in_data[240],
                             in_data[260]};
    
    wire lut_2245_out = lut_2245_table[lut_2245_select];
    
    generate
    if ( USE_REG ) begin : ff_2245
        reg   lut_2245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2245_ff <= lut_2245_out;
            end
        end
        
        assign out_data[2245] = lut_2245_ff;
    end
    else begin : no_ff_2245
        assign out_data[2245] = lut_2245_out;
    end
    endgenerate
    
    
    
    // LUT : 2246
    wire [63:0] lut_2246_table = 64'b0000000000000000000000000001000100000000010101110101010111111111;
    wire [5:0] lut_2246_select = {
                             in_data[513],
                             in_data[407],
                             in_data[485],
                             in_data[532],
                             in_data[55],
                             in_data[211]};
    
    wire lut_2246_out = lut_2246_table[lut_2246_select];
    
    generate
    if ( USE_REG ) begin : ff_2246
        reg   lut_2246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2246_ff <= lut_2246_out;
            end
        end
        
        assign out_data[2246] = lut_2246_ff;
    end
    else begin : no_ff_2246
        assign out_data[2246] = lut_2246_out;
    end
    endgenerate
    
    
    
    // LUT : 2247
    wire [63:0] lut_2247_table = 64'b1110111010001000110011001000100011111111101110111101111111001100;
    wire [5:0] lut_2247_select = {
                             in_data[273],
                             in_data[182],
                             in_data[498],
                             in_data[193],
                             in_data[237],
                             in_data[543]};
    
    wire lut_2247_out = lut_2247_table[lut_2247_select];
    
    generate
    if ( USE_REG ) begin : ff_2247
        reg   lut_2247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2247_ff <= lut_2247_out;
            end
        end
        
        assign out_data[2247] = lut_2247_ff;
    end
    else begin : no_ff_2247
        assign out_data[2247] = lut_2247_out;
    end
    endgenerate
    
    
    
    // LUT : 2248
    wire [63:0] lut_2248_table = 64'b0000000000000000000000000000000000110000101100001111000011110000;
    wire [5:0] lut_2248_select = {
                             in_data[555],
                             in_data[506],
                             in_data[251],
                             in_data[408],
                             in_data[774],
                             in_data[61]};
    
    wire lut_2248_out = lut_2248_table[lut_2248_select];
    
    generate
    if ( USE_REG ) begin : ff_2248
        reg   lut_2248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2248_ff <= lut_2248_out;
            end
        end
        
        assign out_data[2248] = lut_2248_ff;
    end
    else begin : no_ff_2248
        assign out_data[2248] = lut_2248_out;
    end
    endgenerate
    
    
    
    // LUT : 2249
    wire [63:0] lut_2249_table = 64'b1111111101011111111111110101010110110010000000001011000000000000;
    wire [5:0] lut_2249_select = {
                             in_data[373],
                             in_data[520],
                             in_data[637],
                             in_data[286],
                             in_data[60],
                             in_data[552]};
    
    wire lut_2249_out = lut_2249_table[lut_2249_select];
    
    generate
    if ( USE_REG ) begin : ff_2249
        reg   lut_2249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2249_ff <= lut_2249_out;
            end
        end
        
        assign out_data[2249] = lut_2249_ff;
    end
    else begin : no_ff_2249
        assign out_data[2249] = lut_2249_out;
    end
    endgenerate
    
    
    
    // LUT : 2250
    wire [63:0] lut_2250_table = 64'b1111111111111111111111011111110111011100110111001111110011011100;
    wire [5:0] lut_2250_select = {
                             in_data[103],
                             in_data[781],
                             in_data[476],
                             in_data[450],
                             in_data[581],
                             in_data[257]};
    
    wire lut_2250_out = lut_2250_table[lut_2250_select];
    
    generate
    if ( USE_REG ) begin : ff_2250
        reg   lut_2250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2250_ff <= lut_2250_out;
            end
        end
        
        assign out_data[2250] = lut_2250_ff;
    end
    else begin : no_ff_2250
        assign out_data[2250] = lut_2250_out;
    end
    endgenerate
    
    
    
    // LUT : 2251
    wire [63:0] lut_2251_table = 64'b1100111111001111110011111100111111001111110011111100111111001111;
    wire [5:0] lut_2251_select = {
                             in_data[588],
                             in_data[47],
                             in_data[669],
                             in_data[216],
                             in_data[472],
                             in_data[4]};
    
    wire lut_2251_out = lut_2251_table[lut_2251_select];
    
    generate
    if ( USE_REG ) begin : ff_2251
        reg   lut_2251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2251_ff <= lut_2251_out;
            end
        end
        
        assign out_data[2251] = lut_2251_ff;
    end
    else begin : no_ff_2251
        assign out_data[2251] = lut_2251_out;
    end
    endgenerate
    
    
    
    // LUT : 2252
    wire [63:0] lut_2252_table = 64'b0101010101110101010100010011001101010101011101010101000100110011;
    wire [5:0] lut_2252_select = {
                             in_data[36],
                             in_data[147],
                             in_data[179],
                             in_data[539],
                             in_data[298],
                             in_data[322]};
    
    wire lut_2252_out = lut_2252_table[lut_2252_select];
    
    generate
    if ( USE_REG ) begin : ff_2252
        reg   lut_2252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2252_ff <= lut_2252_out;
            end
        end
        
        assign out_data[2252] = lut_2252_ff;
    end
    else begin : no_ff_2252
        assign out_data[2252] = lut_2252_out;
    end
    endgenerate
    
    
    
    // LUT : 2253
    wire [63:0] lut_2253_table = 64'b1111111111001111110011001100110011111111110111111101110011001100;
    wire [5:0] lut_2253_select = {
                             in_data[736],
                             in_data[161],
                             in_data[136],
                             in_data[461],
                             in_data[688],
                             in_data[199]};
    
    wire lut_2253_out = lut_2253_table[lut_2253_select];
    
    generate
    if ( USE_REG ) begin : ff_2253
        reg   lut_2253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2253_ff <= lut_2253_out;
            end
        end
        
        assign out_data[2253] = lut_2253_ff;
    end
    else begin : no_ff_2253
        assign out_data[2253] = lut_2253_out;
    end
    endgenerate
    
    
    
    // LUT : 2254
    wire [63:0] lut_2254_table = 64'b1111101011110000111110101111000011111111111111111111111111110111;
    wire [5:0] lut_2254_select = {
                             in_data[236],
                             in_data[167],
                             in_data[650],
                             in_data[716],
                             in_data[42],
                             in_data[540]};
    
    wire lut_2254_out = lut_2254_table[lut_2254_select];
    
    generate
    if ( USE_REG ) begin : ff_2254
        reg   lut_2254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2254_ff <= lut_2254_out;
            end
        end
        
        assign out_data[2254] = lut_2254_ff;
    end
    else begin : no_ff_2254
        assign out_data[2254] = lut_2254_out;
    end
    endgenerate
    
    
    
    // LUT : 2255
    wire [63:0] lut_2255_table = 64'b0000000000000000000000000000000000000000110000000000000011111111;
    wire [5:0] lut_2255_select = {
                             in_data[121],
                             in_data[333],
                             in_data[178],
                             in_data[765],
                             in_data[717],
                             in_data[783]};
    
    wire lut_2255_out = lut_2255_table[lut_2255_select];
    
    generate
    if ( USE_REG ) begin : ff_2255
        reg   lut_2255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2255_ff <= lut_2255_out;
            end
        end
        
        assign out_data[2255] = lut_2255_ff;
    end
    else begin : no_ff_2255
        assign out_data[2255] = lut_2255_out;
    end
    endgenerate
    
    
    
    // LUT : 2256
    wire [63:0] lut_2256_table = 64'b0000111100000011000011110000111100000000000000000000000000000000;
    wire [5:0] lut_2256_select = {
                             in_data[494],
                             in_data[705],
                             in_data[283],
                             in_data[230],
                             in_data[361],
                             in_data[25]};
    
    wire lut_2256_out = lut_2256_table[lut_2256_select];
    
    generate
    if ( USE_REG ) begin : ff_2256
        reg   lut_2256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2256_ff <= lut_2256_out;
            end
        end
        
        assign out_data[2256] = lut_2256_ff;
    end
    else begin : no_ff_2256
        assign out_data[2256] = lut_2256_out;
    end
    endgenerate
    
    
    
    // LUT : 2257
    wire [63:0] lut_2257_table = 64'b0000000011011100110011001111110011110100110111001111110111011100;
    wire [5:0] lut_2257_select = {
                             in_data[410],
                             in_data[679],
                             in_data[542],
                             in_data[603],
                             in_data[605],
                             in_data[111]};
    
    wire lut_2257_out = lut_2257_table[lut_2257_select];
    
    generate
    if ( USE_REG ) begin : ff_2257
        reg   lut_2257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2257_ff <= lut_2257_out;
            end
        end
        
        assign out_data[2257] = lut_2257_ff;
    end
    else begin : no_ff_2257
        assign out_data[2257] = lut_2257_out;
    end
    endgenerate
    
    
    
    // LUT : 2258
    wire [63:0] lut_2258_table = 64'b1111010011110100111111111111111111110101111100000111000011110000;
    wire [5:0] lut_2258_select = {
                             in_data[526],
                             in_data[442],
                             in_data[26],
                             in_data[624],
                             in_data[757],
                             in_data[722]};
    
    wire lut_2258_out = lut_2258_table[lut_2258_select];
    
    generate
    if ( USE_REG ) begin : ff_2258
        reg   lut_2258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2258_ff <= lut_2258_out;
            end
        end
        
        assign out_data[2258] = lut_2258_ff;
    end
    else begin : no_ff_2258
        assign out_data[2258] = lut_2258_out;
    end
    endgenerate
    
    
    
    // LUT : 2259
    wire [63:0] lut_2259_table = 64'b0101111101000101010101010000010101011111010101010101010100000101;
    wire [5:0] lut_2259_select = {
                             in_data[54],
                             in_data[769],
                             in_data[665],
                             in_data[319],
                             in_data[778],
                             in_data[348]};
    
    wire lut_2259_out = lut_2259_table[lut_2259_select];
    
    generate
    if ( USE_REG ) begin : ff_2259
        reg   lut_2259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2259_ff <= lut_2259_out;
            end
        end
        
        assign out_data[2259] = lut_2259_ff;
    end
    else begin : no_ff_2259
        assign out_data[2259] = lut_2259_out;
    end
    endgenerate
    
    
    
    // LUT : 2260
    wire [63:0] lut_2260_table = 64'b1111111111111111101010101111111100000000111101111010000011111111;
    wire [5:0] lut_2260_select = {
                             in_data[432],
                             in_data[204],
                             in_data[428],
                             in_data[194],
                             in_data[755],
                             in_data[247]};
    
    wire lut_2260_out = lut_2260_table[lut_2260_select];
    
    generate
    if ( USE_REG ) begin : ff_2260
        reg   lut_2260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2260_ff <= lut_2260_out;
            end
        end
        
        assign out_data[2260] = lut_2260_ff;
    end
    else begin : no_ff_2260
        assign out_data[2260] = lut_2260_out;
    end
    endgenerate
    
    
    
    // LUT : 2261
    wire [63:0] lut_2261_table = 64'b1111111100000000000100110000000011111111001000001111001111110010;
    wire [5:0] lut_2261_select = {
                             in_data[403],
                             in_data[242],
                             in_data[354],
                             in_data[122],
                             in_data[583],
                             in_data[479]};
    
    wire lut_2261_out = lut_2261_table[lut_2261_select];
    
    generate
    if ( USE_REG ) begin : ff_2261
        reg   lut_2261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2261_ff <= lut_2261_out;
            end
        end
        
        assign out_data[2261] = lut_2261_ff;
    end
    else begin : no_ff_2261
        assign out_data[2261] = lut_2261_out;
    end
    endgenerate
    
    
    
    // LUT : 2262
    wire [63:0] lut_2262_table = 64'b0001111100011111000011010000110000011111000111110000110100001100;
    wire [5:0] lut_2262_select = {
                             in_data[762],
                             in_data[490],
                             in_data[773],
                             in_data[372],
                             in_data[515],
                             in_data[154]};
    
    wire lut_2262_out = lut_2262_table[lut_2262_select];
    
    generate
    if ( USE_REG ) begin : ff_2262
        reg   lut_2262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2262_ff <= lut_2262_out;
            end
        end
        
        assign out_data[2262] = lut_2262_ff;
    end
    else begin : no_ff_2262
        assign out_data[2262] = lut_2262_out;
    end
    endgenerate
    
    
    
    // LUT : 2263
    wire [63:0] lut_2263_table = 64'b1110111011001100110011001100000011111111111111111111111111111100;
    wire [5:0] lut_2263_select = {
                             in_data[710],
                             in_data[620],
                             in_data[451],
                             in_data[205],
                             in_data[95],
                             in_data[729]};
    
    wire lut_2263_out = lut_2263_table[lut_2263_select];
    
    generate
    if ( USE_REG ) begin : ff_2263
        reg   lut_2263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2263_ff <= lut_2263_out;
            end
        end
        
        assign out_data[2263] = lut_2263_ff;
    end
    else begin : no_ff_2263
        assign out_data[2263] = lut_2263_out;
    end
    endgenerate
    
    
    
    // LUT : 2264
    wire [63:0] lut_2264_table = 64'b0011001000110011001100110011001100110011001100110011001100110011;
    wire [5:0] lut_2264_select = {
                             in_data[52],
                             in_data[336],
                             in_data[686],
                             in_data[172],
                             in_data[523],
                             in_data[768]};
    
    wire lut_2264_out = lut_2264_table[lut_2264_select];
    
    generate
    if ( USE_REG ) begin : ff_2264
        reg   lut_2264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2264_ff <= lut_2264_out;
            end
        end
        
        assign out_data[2264] = lut_2264_ff;
    end
    else begin : no_ff_2264
        assign out_data[2264] = lut_2264_out;
    end
    endgenerate
    
    
    
    // LUT : 2265
    wire [63:0] lut_2265_table = 64'b1100111111001111110011111100111111001111110011111100111111001111;
    wire [5:0] lut_2265_select = {
                             in_data[75],
                             in_data[621],
                             in_data[116],
                             in_data[215],
                             in_data[203],
                             in_data[82]};
    
    wire lut_2265_out = lut_2265_table[lut_2265_select];
    
    generate
    if ( USE_REG ) begin : ff_2265
        reg   lut_2265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2265_ff <= lut_2265_out;
            end
        end
        
        assign out_data[2265] = lut_2265_ff;
    end
    else begin : no_ff_2265
        assign out_data[2265] = lut_2265_out;
    end
    endgenerate
    
    
    
    // LUT : 2266
    wire [63:0] lut_2266_table = 64'b1111111100000010111111110000101010101111000011111010111100001111;
    wire [5:0] lut_2266_select = {
                             in_data[409],
                             in_data[644],
                             in_data[609],
                             in_data[411],
                             in_data[11],
                             in_data[208]};
    
    wire lut_2266_out = lut_2266_table[lut_2266_select];
    
    generate
    if ( USE_REG ) begin : ff_2266
        reg   lut_2266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2266_ff <= lut_2266_out;
            end
        end
        
        assign out_data[2266] = lut_2266_ff;
    end
    else begin : no_ff_2266
        assign out_data[2266] = lut_2266_out;
    end
    endgenerate
    
    
    
    // LUT : 2267
    wire [63:0] lut_2267_table = 64'b1111000011110000100010101000101011110000111100001000101010001110;
    wire [5:0] lut_2267_select = {
                             in_data[50],
                             in_data[345],
                             in_data[779],
                             in_data[292],
                             in_data[239],
                             in_data[234]};
    
    wire lut_2267_out = lut_2267_table[lut_2267_select];
    
    generate
    if ( USE_REG ) begin : ff_2267
        reg   lut_2267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2267_ff <= lut_2267_out;
            end
        end
        
        assign out_data[2267] = lut_2267_ff;
    end
    else begin : no_ff_2267
        assign out_data[2267] = lut_2267_out;
    end
    endgenerate
    
    
    
    // LUT : 2268
    wire [63:0] lut_2268_table = 64'b0000000000000000000000000000000011111111111111111111111111111111;
    wire [5:0] lut_2268_select = {
                             in_data[525],
                             in_data[751],
                             in_data[465],
                             in_data[57],
                             in_data[105],
                             in_data[113]};
    
    wire lut_2268_out = lut_2268_table[lut_2268_select];
    
    generate
    if ( USE_REG ) begin : ff_2268
        reg   lut_2268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2268_ff <= lut_2268_out;
            end
        end
        
        assign out_data[2268] = lut_2268_ff;
    end
    else begin : no_ff_2268
        assign out_data[2268] = lut_2268_out;
    end
    endgenerate
    
    
    
    // LUT : 2269
    wire [63:0] lut_2269_table = 64'b0000100010001100000010001000110000000100010011000000110001001100;
    wire [5:0] lut_2269_select = {
                             in_data[404],
                             in_data[363],
                             in_data[508],
                             in_data[285],
                             in_data[238],
                             in_data[715]};
    
    wire lut_2269_out = lut_2269_table[lut_2269_select];
    
    generate
    if ( USE_REG ) begin : ff_2269
        reg   lut_2269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2269_ff <= lut_2269_out;
            end
        end
        
        assign out_data[2269] = lut_2269_ff;
    end
    else begin : no_ff_2269
        assign out_data[2269] = lut_2269_out;
    end
    endgenerate
    
    
    
    // LUT : 2270
    wire [63:0] lut_2270_table = 64'b1111111111111111111111111111111111111111101010101111101110101010;
    wire [5:0] lut_2270_select = {
                             in_data[426],
                             in_data[533],
                             in_data[129],
                             in_data[2],
                             in_data[88],
                             in_data[664]};
    
    wire lut_2270_out = lut_2270_table[lut_2270_select];
    
    generate
    if ( USE_REG ) begin : ff_2270
        reg   lut_2270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2270_ff <= lut_2270_out;
            end
        end
        
        assign out_data[2270] = lut_2270_ff;
    end
    else begin : no_ff_2270
        assign out_data[2270] = lut_2270_out;
    end
    endgenerate
    
    
    
    // LUT : 2271
    wire [63:0] lut_2271_table = 64'b1111110100000000111111111111111111001100000000001111111111111111;
    wire [5:0] lut_2271_select = {
                             in_data[606],
                             in_data[437],
                             in_data[486],
                             in_data[394],
                             in_data[395],
                             in_data[562]};
    
    wire lut_2271_out = lut_2271_table[lut_2271_select];
    
    generate
    if ( USE_REG ) begin : ff_2271
        reg   lut_2271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2271_ff <= lut_2271_out;
            end
        end
        
        assign out_data[2271] = lut_2271_ff;
    end
    else begin : no_ff_2271
        assign out_data[2271] = lut_2271_out;
    end
    endgenerate
    
    
    
    // LUT : 2272
    wire [63:0] lut_2272_table = 64'b0101010100000000010101010000000001010101000000000101010100000000;
    wire [5:0] lut_2272_select = {
                             in_data[616],
                             in_data[500],
                             in_data[320],
                             in_data[94],
                             in_data[760],
                             in_data[415]};
    
    wire lut_2272_out = lut_2272_table[lut_2272_select];
    
    generate
    if ( USE_REG ) begin : ff_2272
        reg   lut_2272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2272_ff <= lut_2272_out;
            end
        end
        
        assign out_data[2272] = lut_2272_ff;
    end
    else begin : no_ff_2272
        assign out_data[2272] = lut_2272_out;
    end
    endgenerate
    
    
    
    // LUT : 2273
    wire [63:0] lut_2273_table = 64'b0000000000000000000000000000000011111111000100111111111111111111;
    wire [5:0] lut_2273_select = {
                             in_data[315],
                             in_data[402],
                             in_data[590],
                             in_data[22],
                             in_data[86],
                             in_data[560]};
    
    wire lut_2273_out = lut_2273_table[lut_2273_select];
    
    generate
    if ( USE_REG ) begin : ff_2273
        reg   lut_2273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2273_ff <= lut_2273_out;
            end
        end
        
        assign out_data[2273] = lut_2273_ff;
    end
    else begin : no_ff_2273
        assign out_data[2273] = lut_2273_out;
    end
    endgenerate
    
    
    
    // LUT : 2274
    wire [63:0] lut_2274_table = 64'b0000000000000000000100011111101100000000000000000011001111111011;
    wire [5:0] lut_2274_select = {
                             in_data[446],
                             in_data[436],
                             in_data[126],
                             in_data[683],
                             in_data[427],
                             in_data[499]};
    
    wire lut_2274_out = lut_2274_table[lut_2274_select];
    
    generate
    if ( USE_REG ) begin : ff_2274
        reg   lut_2274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2274_ff <= lut_2274_out;
            end
        end
        
        assign out_data[2274] = lut_2274_ff;
    end
    else begin : no_ff_2274
        assign out_data[2274] = lut_2274_out;
    end
    endgenerate
    
    
    
    // LUT : 2275
    wire [63:0] lut_2275_table = 64'b1111111111111111111111111111111111111111010100001111111101010000;
    wire [5:0] lut_2275_select = {
                             in_data[638],
                             in_data[613],
                             in_data[304],
                             in_data[346],
                             in_data[48],
                             in_data[338]};
    
    wire lut_2275_out = lut_2275_table[lut_2275_select];
    
    generate
    if ( USE_REG ) begin : ff_2275
        reg   lut_2275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2275_ff <= lut_2275_out;
            end
        end
        
        assign out_data[2275] = lut_2275_ff;
    end
    else begin : no_ff_2275
        assign out_data[2275] = lut_2275_out;
    end
    endgenerate
    
    
    
    // LUT : 2276
    wire [63:0] lut_2276_table = 64'b1111111100000000111111110000000011111111000000001111111100000000;
    wire [5:0] lut_2276_select = {
                             in_data[693],
                             in_data[584],
                             in_data[470],
                             in_data[46],
                             in_data[599],
                             in_data[720]};
    
    wire lut_2276_out = lut_2276_table[lut_2276_select];
    
    generate
    if ( USE_REG ) begin : ff_2276
        reg   lut_2276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2276_ff <= lut_2276_out;
            end
        end
        
        assign out_data[2276] = lut_2276_ff;
    end
    else begin : no_ff_2276
        assign out_data[2276] = lut_2276_out;
    end
    endgenerate
    
    
    
    // LUT : 2277
    wire [63:0] lut_2277_table = 64'b0000000000000000000000000000000000100010111011100010001010101010;
    wire [5:0] lut_2277_select = {
                             in_data[567],
                             in_data[6],
                             in_data[537],
                             in_data[780],
                             in_data[189],
                             in_data[430]};
    
    wire lut_2277_out = lut_2277_table[lut_2277_select];
    
    generate
    if ( USE_REG ) begin : ff_2277
        reg   lut_2277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2277_ff <= lut_2277_out;
            end
        end
        
        assign out_data[2277] = lut_2277_ff;
    end
    else begin : no_ff_2277
        assign out_data[2277] = lut_2277_out;
    end
    endgenerate
    
    
    
    // LUT : 2278
    wire [63:0] lut_2278_table = 64'b0010000000100000001000001011000010110010101100111011001010110010;
    wire [5:0] lut_2278_select = {
                             in_data[608],
                             in_data[389],
                             in_data[702],
                             in_data[625],
                             in_data[400],
                             in_data[356]};
    
    wire lut_2278_out = lut_2278_table[lut_2278_select];
    
    generate
    if ( USE_REG ) begin : ff_2278
        reg   lut_2278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2278_ff <= lut_2278_out;
            end
        end
        
        assign out_data[2278] = lut_2278_ff;
    end
    else begin : no_ff_2278
        assign out_data[2278] = lut_2278_out;
    end
    endgenerate
    
    
    
    // LUT : 2279
    wire [63:0] lut_2279_table = 64'b0101000011111111010100000111011101010000111111110000000001110111;
    wire [5:0] lut_2279_select = {
                             in_data[393],
                             in_data[544],
                             in_data[351],
                             in_data[149],
                             in_data[595],
                             in_data[382]};
    
    wire lut_2279_out = lut_2279_table[lut_2279_select];
    
    generate
    if ( USE_REG ) begin : ff_2279
        reg   lut_2279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2279_ff <= lut_2279_out;
            end
        end
        
        assign out_data[2279] = lut_2279_ff;
    end
    else begin : no_ff_2279
        assign out_data[2279] = lut_2279_out;
    end
    endgenerate
    
    
    
    // LUT : 2280
    wire [63:0] lut_2280_table = 64'b1111111111111111111111001111110011111111111111111111110011111100;
    wire [5:0] lut_2280_select = {
                             in_data[67],
                             in_data[268],
                             in_data[337],
                             in_data[714],
                             in_data[737],
                             in_data[140]};
    
    wire lut_2280_out = lut_2280_table[lut_2280_select];
    
    generate
    if ( USE_REG ) begin : ff_2280
        reg   lut_2280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2280_ff <= lut_2280_out;
            end
        end
        
        assign out_data[2280] = lut_2280_ff;
    end
    else begin : no_ff_2280
        assign out_data[2280] = lut_2280_out;
    end
    endgenerate
    
    
    
    // LUT : 2281
    wire [63:0] lut_2281_table = 64'b0000001100110011001100110011000000000011001100000011001100110011;
    wire [5:0] lut_2281_select = {
                             in_data[478],
                             in_data[766],
                             in_data[496],
                             in_data[155],
                             in_data[232],
                             in_data[727]};
    
    wire lut_2281_out = lut_2281_table[lut_2281_select];
    
    generate
    if ( USE_REG ) begin : ff_2281
        reg   lut_2281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2281_ff <= lut_2281_out;
            end
        end
        
        assign out_data[2281] = lut_2281_ff;
    end
    else begin : no_ff_2281
        assign out_data[2281] = lut_2281_out;
    end
    endgenerate
    
    
    
    // LUT : 2282
    wire [63:0] lut_2282_table = 64'b1111000011110000111100000000000011111111111100001111000011110000;
    wire [5:0] lut_2282_select = {
                             in_data[723],
                             in_data[529],
                             in_data[185],
                             in_data[598],
                             in_data[109],
                             in_data[646]};
    
    wire lut_2282_out = lut_2282_table[lut_2282_select];
    
    generate
    if ( USE_REG ) begin : ff_2282
        reg   lut_2282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2282_ff <= lut_2282_out;
            end
        end
        
        assign out_data[2282] = lut_2282_ff;
    end
    else begin : no_ff_2282
        assign out_data[2282] = lut_2282_out;
    end
    endgenerate
    
    
    
    // LUT : 2283
    wire [63:0] lut_2283_table = 64'b0000000001000101010000001100000011100100111101011111010011110100;
    wire [5:0] lut_2283_select = {
                             in_data[213],
                             in_data[433],
                             in_data[711],
                             in_data[548],
                             in_data[740],
                             in_data[150]};
    
    wire lut_2283_out = lut_2283_table[lut_2283_select];
    
    generate
    if ( USE_REG ) begin : ff_2283
        reg   lut_2283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2283_ff <= lut_2283_out;
            end
        end
        
        assign out_data[2283] = lut_2283_ff;
    end
    else begin : no_ff_2283
        assign out_data[2283] = lut_2283_out;
    end
    endgenerate
    
    
    
    // LUT : 2284
    wire [63:0] lut_2284_table = 64'b1111000011111111111100001111000011110000111111111111000011110000;
    wire [5:0] lut_2284_select = {
                             in_data[78],
                             in_data[467],
                             in_data[458],
                             in_data[607],
                             in_data[447],
                             in_data[618]};
    
    wire lut_2284_out = lut_2284_table[lut_2284_select];
    
    generate
    if ( USE_REG ) begin : ff_2284
        reg   lut_2284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2284_ff <= lut_2284_out;
            end
        end
        
        assign out_data[2284] = lut_2284_ff;
    end
    else begin : no_ff_2284
        assign out_data[2284] = lut_2284_out;
    end
    endgenerate
    
    
    
    // LUT : 2285
    wire [63:0] lut_2285_table = 64'b0101010111110101010101011111010101010101010101010101010101010101;
    wire [5:0] lut_2285_select = {
                             in_data[687],
                             in_data[501],
                             in_data[680],
                             in_data[739],
                             in_data[170],
                             in_data[511]};
    
    wire lut_2285_out = lut_2285_table[lut_2285_select];
    
    generate
    if ( USE_REG ) begin : ff_2285
        reg   lut_2285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2285_ff <= lut_2285_out;
            end
        end
        
        assign out_data[2285] = lut_2285_ff;
    end
    else begin : no_ff_2285
        assign out_data[2285] = lut_2285_out;
    end
    endgenerate
    
    
    
    // LUT : 2286
    wire [63:0] lut_2286_table = 64'b1010101010101010001000100010001011111011111110111011101110111011;
    wire [5:0] lut_2286_select = {
                             in_data[184],
                             in_data[66],
                             in_data[114],
                             in_data[37],
                             in_data[719],
                             in_data[651]};
    
    wire lut_2286_out = lut_2286_table[lut_2286_select];
    
    generate
    if ( USE_REG ) begin : ff_2286
        reg   lut_2286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2286_ff <= lut_2286_out;
            end
        end
        
        assign out_data[2286] = lut_2286_ff;
    end
    else begin : no_ff_2286
        assign out_data[2286] = lut_2286_out;
    end
    endgenerate
    
    
    
    // LUT : 2287
    wire [63:0] lut_2287_table = 64'b1111111111111111111111111111111101011111010100001111101011111010;
    wire [5:0] lut_2287_select = {
                             in_data[340],
                             in_data[656],
                             in_data[93],
                             in_data[681],
                             in_data[51],
                             in_data[575]};
    
    wire lut_2287_out = lut_2287_table[lut_2287_select];
    
    generate
    if ( USE_REG ) begin : ff_2287
        reg   lut_2287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2287_ff <= lut_2287_out;
            end
        end
        
        assign out_data[2287] = lut_2287_ff;
    end
    else begin : no_ff_2287
        assign out_data[2287] = lut_2287_out;
    end
    endgenerate
    
    
    
    // LUT : 2288
    wire [63:0] lut_2288_table = 64'b0011000000110000000111110000111100100000001000000000111100011111;
    wire [5:0] lut_2288_select = {
                             in_data[38],
                             in_data[438],
                             in_data[39],
                             in_data[375],
                             in_data[471],
                             in_data[325]};
    
    wire lut_2288_out = lut_2288_table[lut_2288_select];
    
    generate
    if ( USE_REG ) begin : ff_2288
        reg   lut_2288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2288_ff <= lut_2288_out;
            end
        end
        
        assign out_data[2288] = lut_2288_ff;
    end
    else begin : no_ff_2288
        assign out_data[2288] = lut_2288_out;
    end
    endgenerate
    
    
    
    // LUT : 2289
    wire [63:0] lut_2289_table = 64'b1010101010101010101010101010101010101010101010101010111010101010;
    wire [5:0] lut_2289_select = {
                             in_data[288],
                             in_data[753],
                             in_data[612],
                             in_data[8],
                             in_data[640],
                             in_data[187]};
    
    wire lut_2289_out = lut_2289_table[lut_2289_select];
    
    generate
    if ( USE_REG ) begin : ff_2289
        reg   lut_2289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2289_ff <= lut_2289_out;
            end
        end
        
        assign out_data[2289] = lut_2289_ff;
    end
    else begin : no_ff_2289
        assign out_data[2289] = lut_2289_out;
    end
    endgenerate
    
    
    
    // LUT : 2290
    wire [63:0] lut_2290_table = 64'b1111111111111111111110001111100011111111111111111111101011111010;
    wire [5:0] lut_2290_select = {
                             in_data[138],
                             in_data[294],
                             in_data[713],
                             in_data[227],
                             in_data[502],
                             in_data[648]};
    
    wire lut_2290_out = lut_2290_table[lut_2290_select];
    
    generate
    if ( USE_REG ) begin : ff_2290
        reg   lut_2290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2290_ff <= lut_2290_out;
            end
        end
        
        assign out_data[2290] = lut_2290_ff;
    end
    else begin : no_ff_2290
        assign out_data[2290] = lut_2290_out;
    end
    endgenerate
    
    
    
    // LUT : 2291
    wire [63:0] lut_2291_table = 64'b0000111110101111000000000000000011111111111111110000100000000000;
    wire [5:0] lut_2291_select = {
                             in_data[586],
                             in_data[601],
                             in_data[704],
                             in_data[159],
                             in_data[10],
                             in_data[734]};
    
    wire lut_2291_out = lut_2291_table[lut_2291_select];
    
    generate
    if ( USE_REG ) begin : ff_2291
        reg   lut_2291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2291_ff <= lut_2291_out;
            end
        end
        
        assign out_data[2291] = lut_2291_ff;
    end
    else begin : no_ff_2291
        assign out_data[2291] = lut_2291_out;
    end
    endgenerate
    
    
    
    // LUT : 2292
    wire [63:0] lut_2292_table = 64'b0101011111111111000000000000000011010111111111110000000000000000;
    wire [5:0] lut_2292_select = {
                             in_data[764],
                             in_data[297],
                             in_data[464],
                             in_data[770],
                             in_data[198],
                             in_data[259]};
    
    wire lut_2292_out = lut_2292_table[lut_2292_select];
    
    generate
    if ( USE_REG ) begin : ff_2292
        reg   lut_2292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2292_ff <= lut_2292_out;
            end
        end
        
        assign out_data[2292] = lut_2292_ff;
    end
    else begin : no_ff_2292
        assign out_data[2292] = lut_2292_out;
    end
    endgenerate
    
    
    
    // LUT : 2293
    wire [63:0] lut_2293_table = 64'b1111111111111110111111111111111011111111111111101111111111111110;
    wire [5:0] lut_2293_select = {
                             in_data[699],
                             in_data[27],
                             in_data[691],
                             in_data[148],
                             in_data[480],
                             in_data[90]};
    
    wire lut_2293_out = lut_2293_table[lut_2293_select];
    
    generate
    if ( USE_REG ) begin : ff_2293
        reg   lut_2293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2293_ff <= lut_2293_out;
            end
        end
        
        assign out_data[2293] = lut_2293_ff;
    end
    else begin : no_ff_2293
        assign out_data[2293] = lut_2293_out;
    end
    endgenerate
    
    
    
    // LUT : 2294
    wire [63:0] lut_2294_table = 64'b1111111011111111000000000000000011001100111111111100100011001100;
    wire [5:0] lut_2294_select = {
                             in_data[130],
                             in_data[128],
                             in_data[663],
                             in_data[761],
                             in_data[291],
                             in_data[561]};
    
    wire lut_2294_out = lut_2294_table[lut_2294_select];
    
    generate
    if ( USE_REG ) begin : ff_2294
        reg   lut_2294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2294_ff <= lut_2294_out;
            end
        end
        
        assign out_data[2294] = lut_2294_ff;
    end
    else begin : no_ff_2294
        assign out_data[2294] = lut_2294_out;
    end
    endgenerate
    
    
    
    // LUT : 2295
    wire [63:0] lut_2295_table = 64'b1111001111111011111110111111111111110011111100111111001111110011;
    wire [5:0] lut_2295_select = {
                             in_data[706],
                             in_data[397],
                             in_data[310],
                             in_data[173],
                             in_data[514],
                             in_data[23]};
    
    wire lut_2295_out = lut_2295_table[lut_2295_select];
    
    generate
    if ( USE_REG ) begin : ff_2295
        reg   lut_2295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2295_ff <= lut_2295_out;
            end
        end
        
        assign out_data[2295] = lut_2295_ff;
    end
    else begin : no_ff_2295
        assign out_data[2295] = lut_2295_out;
    end
    endgenerate
    
    
    
    // LUT : 2296
    wire [63:0] lut_2296_table = 64'b0000000000000000000000000000000000000000000000000000001100110011;
    wire [5:0] lut_2296_select = {
                             in_data[70],
                             in_data[399],
                             in_data[572],
                             in_data[682],
                             in_data[398],
                             in_data[422]};
    
    wire lut_2296_out = lut_2296_table[lut_2296_select];
    
    generate
    if ( USE_REG ) begin : ff_2296
        reg   lut_2296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2296_ff <= lut_2296_out;
            end
        end
        
        assign out_data[2296] = lut_2296_ff;
    end
    else begin : no_ff_2296
        assign out_data[2296] = lut_2296_out;
    end
    endgenerate
    
    
    
    // LUT : 2297
    wire [63:0] lut_2297_table = 64'b1111111111111111000000001010000011110001101010101111000110100000;
    wire [5:0] lut_2297_select = {
                             in_data[132],
                             in_data[271],
                             in_data[386],
                             in_data[295],
                             in_data[668],
                             in_data[212]};
    
    wire lut_2297_out = lut_2297_table[lut_2297_select];
    
    generate
    if ( USE_REG ) begin : ff_2297
        reg   lut_2297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2297_ff <= lut_2297_out;
            end
        end
        
        assign out_data[2297] = lut_2297_ff;
    end
    else begin : no_ff_2297
        assign out_data[2297] = lut_2297_out;
    end
    endgenerate
    
    
    
    // LUT : 2298
    wire [63:0] lut_2298_table = 64'b1111110011111100111111111111111100110000001100000011000000110000;
    wire [5:0] lut_2298_select = {
                             in_data[347],
                             in_data[96],
                             in_data[392],
                             in_data[463],
                             in_data[412],
                             in_data[254]};
    
    wire lut_2298_out = lut_2298_table[lut_2298_select];
    
    generate
    if ( USE_REG ) begin : ff_2298
        reg   lut_2298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2298_ff <= lut_2298_out;
            end
        end
        
        assign out_data[2298] = lut_2298_ff;
    end
    else begin : no_ff_2298
        assign out_data[2298] = lut_2298_out;
    end
    endgenerate
    
    
    
    // LUT : 2299
    wire [63:0] lut_2299_table = 64'b0000010000000000000011110000000000001111000000000000111100000101;
    wire [5:0] lut_2299_select = {
                             in_data[225],
                             in_data[107],
                             in_data[674],
                             in_data[250],
                             in_data[558],
                             in_data[521]};
    
    wire lut_2299_out = lut_2299_table[lut_2299_select];
    
    generate
    if ( USE_REG ) begin : ff_2299
        reg   lut_2299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2299_ff <= lut_2299_out;
            end
        end
        
        assign out_data[2299] = lut_2299_ff;
    end
    else begin : no_ff_2299
        assign out_data[2299] = lut_2299_out;
    end
    endgenerate
    
    
    
    // LUT : 2300
    wire [63:0] lut_2300_table = 64'b0111010101010101010101010101010101010101000101010101010100010001;
    wire [5:0] lut_2300_select = {
                             in_data[164],
                             in_data[137],
                             in_data[49],
                             in_data[308],
                             in_data[371],
                             in_data[229]};
    
    wire lut_2300_out = lut_2300_table[lut_2300_select];
    
    generate
    if ( USE_REG ) begin : ff_2300
        reg   lut_2300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2300_ff <= lut_2300_out;
            end
        end
        
        assign out_data[2300] = lut_2300_ff;
    end
    else begin : no_ff_2300
        assign out_data[2300] = lut_2300_out;
    end
    endgenerate
    
    
    
    // LUT : 2301
    wire [63:0] lut_2301_table = 64'b0000000011111111000000000010001010101010111111111010101010101010;
    wire [5:0] lut_2301_select = {
                             in_data[72],
                             in_data[709],
                             in_data[602],
                             in_data[45],
                             in_data[334],
                             in_data[455]};
    
    wire lut_2301_out = lut_2301_table[lut_2301_select];
    
    generate
    if ( USE_REG ) begin : ff_2301
        reg   lut_2301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2301_ff <= lut_2301_out;
            end
        end
        
        assign out_data[2301] = lut_2301_ff;
    end
    else begin : no_ff_2301
        assign out_data[2301] = lut_2301_out;
    end
    endgenerate
    
    
    
    // LUT : 2302
    wire [63:0] lut_2302_table = 64'b1111111111111111111111111111111101010101010101010000000000000000;
    wire [5:0] lut_2302_select = {
                             in_data[443],
                             in_data[547],
                             in_data[83],
                             in_data[307],
                             in_data[366],
                             in_data[658]};
    
    wire lut_2302_out = lut_2302_table[lut_2302_select];
    
    generate
    if ( USE_REG ) begin : ff_2302
        reg   lut_2302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2302_ff <= lut_2302_out;
            end
        end
        
        assign out_data[2302] = lut_2302_ff;
    end
    else begin : no_ff_2302
        assign out_data[2302] = lut_2302_out;
    end
    endgenerate
    
    
    
    // LUT : 2303
    wire [63:0] lut_2303_table = 64'b0000000000000000000000001111111100000000000000000000000011111111;
    wire [5:0] lut_2303_select = {
                             in_data[0],
                             in_data[284],
                             in_data[206],
                             in_data[477],
                             in_data[524],
                             in_data[369]};
    
    wire lut_2303_out = lut_2303_table[lut_2303_select];
    
    generate
    if ( USE_REG ) begin : ff_2303
        reg   lut_2303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2303_ff <= lut_2303_out;
            end
        end
        
        assign out_data[2303] = lut_2303_ff;
    end
    else begin : no_ff_2303
        assign out_data[2303] = lut_2303_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub1
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [       2303:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        383:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub1_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub1_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub1_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [2303:0]  in_data,
            output wire [383:0]  out_data
        );
    
    
    // LUT : 0
    wire [63:0] lut_0_table = 64'b1111110111111111111111000111000000000000000100010001000000010000;
    wire [5:0] lut_0_select = {
                             in_data[111],
                             in_data[1178],
                             in_data[1260],
                             in_data[1485],
                             in_data[302],
                             in_data[531]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [63:0] lut_1_table = 64'b0101111100001110010111010000000001010111000100110111111100010011;
    wire [5:0] lut_1_select = {
                             in_data[1873],
                             in_data[1254],
                             in_data[203],
                             in_data[1074],
                             in_data[1283],
                             in_data[812]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [63:0] lut_2_table = 64'b1111111101010000111111100000000001111010000000101110000000000000;
    wire [5:0] lut_2_select = {
                             in_data[898],
                             in_data[1580],
                             in_data[725],
                             in_data[2242],
                             in_data[1890],
                             in_data[620]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [63:0] lut_3_table = 64'b1000110111001111100011111000111111001110111111111010101110111111;
    wire [5:0] lut_3_select = {
                             in_data[330],
                             in_data[2213],
                             in_data[1728],
                             in_data[1457],
                             in_data[1330],
                             in_data[2135]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [63:0] lut_4_table = 64'b1000100011101100001000100010000010001000110011000010000000001000;
    wire [5:0] lut_4_select = {
                             in_data[932],
                             in_data[1770],
                             in_data[1029],
                             in_data[1777],
                             in_data[742],
                             in_data[2181]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [63:0] lut_5_table = 64'b1101110011101100111111001111110011110000111011001111100011111110;
    wire [5:0] lut_5_select = {
                             in_data[574],
                             in_data[2064],
                             in_data[2047],
                             in_data[193],
                             in_data[1715],
                             in_data[771]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [63:0] lut_6_table = 64'b1111110011000000110000000000000011111110100010001110111010000000;
    wire [5:0] lut_6_select = {
                             in_data[966],
                             in_data[359],
                             in_data[580],
                             in_data[1851],
                             in_data[608],
                             in_data[1629]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [63:0] lut_7_table = 64'b0100000000000000000000000000000011111111010011000100110000000000;
    wire [5:0] lut_7_select = {
                             in_data[1751],
                             in_data[2108],
                             in_data[1566],
                             in_data[1882],
                             in_data[320],
                             in_data[1543]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [63:0] lut_8_table = 64'b1111111111010000011100010100000001110111011110110000001100000000;
    wire [5:0] lut_8_select = {
                             in_data[1182],
                             in_data[101],
                             in_data[2152],
                             in_data[490],
                             in_data[2203],
                             in_data[1913]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [63:0] lut_9_table = 64'b0010000011101000000000001111111000001010010011000000110011001100;
    wire [5:0] lut_9_select = {
                             in_data[1973],
                             in_data[322],
                             in_data[745],
                             in_data[472],
                             in_data[141],
                             in_data[972]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [63:0] lut_10_table = 64'b1111110111111111111111110111111101000000010001001100110001001101;
    wire [5:0] lut_10_select = {
                             in_data[2188],
                             in_data[1726],
                             in_data[252],
                             in_data[522],
                             in_data[2218],
                             in_data[1931]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [63:0] lut_11_table = 64'b0000110000001111000011001100111100000100000011110000110000001111;
    wire [5:0] lut_11_select = {
                             in_data[125],
                             in_data[820],
                             in_data[1671],
                             in_data[1533],
                             in_data[53],
                             in_data[689]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [63:0] lut_12_table = 64'b0000000000001000000111011111111100001000100010000001110111011111;
    wire [5:0] lut_12_select = {
                             in_data[1559],
                             in_data[1968],
                             in_data[340],
                             in_data[602],
                             in_data[171],
                             in_data[789]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [63:0] lut_13_table = 64'b0000001010100010111111111111011101001101000000001101111101000101;
    wire [5:0] lut_13_select = {
                             in_data[1969],
                             in_data[1420],
                             in_data[1215],
                             in_data[1655],
                             in_data[1564],
                             in_data[232]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [63:0] lut_14_table = 64'b1111111111111111111111110001000101110001010100010011001100000000;
    wire [5:0] lut_14_select = {
                             in_data[526],
                             in_data[1201],
                             in_data[1592],
                             in_data[2149],
                             in_data[993],
                             in_data[970]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [63:0] lut_15_table = 64'b1100110111111111111111111111111101001100110111111100110011111111;
    wire [5:0] lut_15_select = {
                             in_data[600],
                             in_data[1199],
                             in_data[267],
                             in_data[1077],
                             in_data[1708],
                             in_data[701]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [63:0] lut_16_table = 64'b0101000000000000011100010001000011110001010101000111001101010001;
    wire [5:0] lut_16_select = {
                             in_data[2157],
                             in_data[116],
                             in_data[2255],
                             in_data[1550],
                             in_data[97],
                             in_data[368]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [63:0] lut_17_table = 64'b0000100000110111000000000001000101001100001111110000000000010101;
    wire [5:0] lut_17_select = {
                             in_data[1695],
                             in_data[1908],
                             in_data[2292],
                             in_data[481],
                             in_data[749],
                             in_data[77]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [63:0] lut_18_table = 64'b1100110000000100111111010000010011001100000000001100110100000100;
    wire [5:0] lut_18_select = {
                             in_data[152],
                             in_data[805],
                             in_data[33],
                             in_data[1088],
                             in_data[374],
                             in_data[1676]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [63:0] lut_19_table = 64'b1100111111011111111111011111111110001000110011101101100011001110;
    wire [5:0] lut_19_select = {
                             in_data[2017],
                             in_data[1611],
                             in_data[1396],
                             in_data[2216],
                             in_data[365],
                             in_data[1509]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [63:0] lut_20_table = 64'b0111011101110111011001100111111001010111000101111111111100111110;
    wire [5:0] lut_20_select = {
                             in_data[64],
                             in_data[852],
                             in_data[436],
                             in_data[427],
                             in_data[172],
                             in_data[393]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [63:0] lut_21_table = 64'b0000000011110111010101111111111101000000010101010100011101001111;
    wire [5:0] lut_21_select = {
                             in_data[2067],
                             in_data[1300],
                             in_data[549],
                             in_data[1731],
                             in_data[1517],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [63:0] lut_22_table = 64'b1110111011111111100010001110110110001000111010111000000010000000;
    wire [5:0] lut_22_select = {
                             in_data[43],
                             in_data[1716],
                             in_data[1553],
                             in_data[628],
                             in_data[1831],
                             in_data[1151]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [63:0] lut_23_table = 64'b0000000000100000000000000000000000000000001100110011000101111111;
    wire [5:0] lut_23_select = {
                             in_data[648],
                             in_data[1583],
                             in_data[924],
                             in_data[1656],
                             in_data[1251],
                             in_data[2286]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [63:0] lut_24_table = 64'b1100000011001000111011001111111010000000100000001100010011101100;
    wire [5:0] lut_24_select = {
                             in_data[511],
                             in_data[1502],
                             in_data[1133],
                             in_data[1597],
                             in_data[1791],
                             in_data[1430]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [63:0] lut_25_table = 64'b0101000101010101000000000000000111110000111101010101000001010000;
    wire [5:0] lut_25_select = {
                             in_data[63],
                             in_data[1764],
                             in_data[1883],
                             in_data[142],
                             in_data[1979],
                             in_data[601]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [63:0] lut_26_table = 64'b0000111101011111000011110000111101011111000011110000111100001110;
    wire [5:0] lut_26_select = {
                             in_data[1775],
                             in_data[1887],
                             in_data[1013],
                             in_data[1977],
                             in_data[179],
                             in_data[131]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [63:0] lut_27_table = 64'b1010101000001111101010101111111100000000000000001010101000001111;
    wire [5:0] lut_27_select = {
                             in_data[1257],
                             in_data[1993],
                             in_data[2165],
                             in_data[223],
                             in_data[521],
                             in_data[432]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [63:0] lut_28_table = 64'b1100101010010000111111111111111000000000000001000000111011111111;
    wire [5:0] lut_28_select = {
                             in_data[1975],
                             in_data[774],
                             in_data[1827],
                             in_data[634],
                             in_data[2],
                             in_data[1282]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [63:0] lut_29_table = 64'b0011111101011111110011110100111101010111000001011111111101001111;
    wire [5:0] lut_29_select = {
                             in_data[2214],
                             in_data[130],
                             in_data[1576],
                             in_data[1495],
                             in_data[1588],
                             in_data[1323]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [63:0] lut_30_table = 64'b0000111100001111111111111111111100001100000001010000011100111111;
    wire [5:0] lut_30_select = {
                             in_data[286],
                             in_data[1248],
                             in_data[415],
                             in_data[2221],
                             in_data[1089],
                             in_data[1510]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [63:0] lut_31_table = 64'b1111100011111010100000001000000011110000111110100011000000110000;
    wire [5:0] lut_31_select = {
                             in_data[228],
                             in_data[1544],
                             in_data[160],
                             in_data[1314],
                             in_data[1350],
                             in_data[649]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [63:0] lut_32_table = 64'b1011111100000000111111110000000000111111000000000000011000000000;
    wire [5:0] lut_32_select = {
                             in_data[1896],
                             in_data[2102],
                             in_data[1538],
                             in_data[2301],
                             in_data[229],
                             in_data[914]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [63:0] lut_33_table = 64'b0000111100001111000010010000000000111111111111110000111100001101;
    wire [5:0] lut_33_select = {
                             in_data[1894],
                             in_data[1466],
                             in_data[318],
                             in_data[1529],
                             in_data[2025],
                             in_data[39]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [63:0] lut_34_table = 64'b0011000000000000101100000000000010111100101111101010100010101010;
    wire [5:0] lut_34_select = {
                             in_data[1234],
                             in_data[1866],
                             in_data[1959],
                             in_data[863],
                             in_data[756],
                             in_data[1563]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [63:0] lut_35_table = 64'b0010111100000000111111110000000011111010000100001111111101110000;
    wire [5:0] lut_35_select = {
                             in_data[190],
                             in_data[2032],
                             in_data[209],
                             in_data[418],
                             in_data[1868],
                             in_data[1720]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [63:0] lut_36_table = 64'b1100000011000000100010101111101001000000110000000000000011111010;
    wire [5:0] lut_36_select = {
                             in_data[1669],
                             in_data[652],
                             in_data[370],
                             in_data[367],
                             in_data[2130],
                             in_data[796]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [63:0] lut_37_table = 64'b1111111100010001010111110000000111111111010100011111111100010111;
    wire [5:0] lut_37_select = {
                             in_data[22],
                             in_data[2230],
                             in_data[1773],
                             in_data[2154],
                             in_data[478],
                             in_data[1456]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [63:0] lut_38_table = 64'b0101000001110111011100111111111100000000010101010111000111111111;
    wire [5:0] lut_38_select = {
                             in_data[818],
                             in_data[851],
                             in_data[886],
                             in_data[1692],
                             in_data[1985],
                             in_data[1127]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [63:0] lut_39_table = 64'b1100110011111111110011011101111101000100110111110101010111011101;
    wire [5:0] lut_39_select = {
                             in_data[1955],
                             in_data[916],
                             in_data[114],
                             in_data[894],
                             in_data[2191],
                             in_data[1369]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [63:0] lut_40_table = 64'b0100010111111111010001001101111100000001111111110000000001000000;
    wire [5:0] lut_40_select = {
                             in_data[364],
                             in_data[173],
                             in_data[326],
                             in_data[603],
                             in_data[1021],
                             in_data[1527]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [63:0] lut_41_table = 64'b1100000011110000100010001000100011110000110000001111111011000000;
    wire [5:0] lut_41_select = {
                             in_data[210],
                             in_data[2070],
                             in_data[473],
                             in_data[913],
                             in_data[956],
                             in_data[1263]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [63:0] lut_42_table = 64'b1111111101110110010001000000000001010100010001000100010001000100;
    wire [5:0] lut_42_select = {
                             in_data[1326],
                             in_data[2200],
                             in_data[887],
                             in_data[1179],
                             in_data[635],
                             in_data[2058]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [63:0] lut_43_table = 64'b0111000011110100111100101111111100000000010000000000000001000100;
    wire [5:0] lut_43_select = {
                             in_data[1382],
                             in_data[1738],
                             in_data[1491],
                             in_data[1754],
                             in_data[1130],
                             in_data[976]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [63:0] lut_44_table = 64'b0000000010101010100010101110111011111111000000001100100010001000;
    wire [5:0] lut_44_select = {
                             in_data[1209],
                             in_data[896],
                             in_data[937],
                             in_data[640],
                             in_data[1208],
                             in_data[1587]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [63:0] lut_45_table = 64'b0000000011011101000001000110111100001101100011110000011100000010;
    wire [5:0] lut_45_select = {
                             in_data[373],
                             in_data[1163],
                             in_data[2048],
                             in_data[1444],
                             in_data[299],
                             in_data[460]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [63:0] lut_46_table = 64'b1100111010001010000010111110111000001000000010000000000010001010;
    wire [5:0] lut_46_select = {
                             in_data[509],
                             in_data[170],
                             in_data[750],
                             in_data[905],
                             in_data[1351],
                             in_data[2298]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [63:0] lut_47_table = 64'b1000101010101010101010110010001010001000000000001010001000000000;
    wire [5:0] lut_47_select = {
                             in_data[297],
                             in_data[1589],
                             in_data[1503],
                             in_data[288],
                             in_data[849],
                             in_data[83]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [63:0] lut_48_table = 64'b0000111100010111111111111111111100000000000000001111111111111011;
    wire [5:0] lut_48_select = {
                             in_data[930],
                             in_data[184],
                             in_data[117],
                             in_data[1183],
                             in_data[2040],
                             in_data[1214]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [63:0] lut_49_table = 64'b0101010101110101000100000111000100110000001100000011000001110000;
    wire [5:0] lut_49_select = {
                             in_data[1750],
                             in_data[1710],
                             in_data[1911],
                             in_data[856],
                             in_data[822],
                             in_data[56]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [63:0] lut_50_table = 64'b0000001000000000111111110000000011001111010001001100111100001100;
    wire [5:0] lut_50_select = {
                             in_data[306],
                             in_data[1621],
                             in_data[1309],
                             in_data[1938],
                             in_data[458],
                             in_data[1749]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [63:0] lut_51_table = 64'b1111000111110101111100001111000011110000111100000011000010110000;
    wire [5:0] lut_51_select = {
                             in_data[1333],
                             in_data[213],
                             in_data[797],
                             in_data[925],
                             in_data[566],
                             in_data[902]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [63:0] lut_52_table = 64'b0001001100011011000000001111111100010011000100010000000011011101;
    wire [5:0] lut_52_select = {
                             in_data[165],
                             in_data[572],
                             in_data[1598],
                             in_data[638],
                             in_data[1943],
                             in_data[423]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [63:0] lut_53_table = 64'b0001111100001111111111111000110100000001000011010101010100000101;
    wire [5:0] lut_53_select = {
                             in_data[7],
                             in_data[667],
                             in_data[1619],
                             in_data[1311],
                             in_data[2302],
                             in_data[895]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [63:0] lut_54_table = 64'b1111111100001111010011110000010011111111010001010101110101000100;
    wire [5:0] lut_54_select = {
                             in_data[1156],
                             in_data[313],
                             in_data[1020],
                             in_data[6],
                             in_data[1229],
                             in_data[2189]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [63:0] lut_55_table = 64'b0000101000000000101000101110000010101010111100101000000011110000;
    wire [5:0] lut_55_select = {
                             in_data[255],
                             in_data[1888],
                             in_data[637],
                             in_data[527],
                             in_data[18],
                             in_data[1272]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [63:0] lut_56_table = 64'b1100110010001100110011001100110011001100111011101100111011001100;
    wire [5:0] lut_56_select = {
                             in_data[2248],
                             in_data[217],
                             in_data[106],
                             in_data[1167],
                             in_data[2099],
                             in_data[757]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [63:0] lut_57_table = 64'b1100010001000000110001000000000011111101111101001100110011000100;
    wire [5:0] lut_57_select = {
                             in_data[726],
                             in_data[146],
                             in_data[1389],
                             in_data[242],
                             in_data[1983],
                             in_data[650]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [63:0] lut_58_table = 64'b0000000010100000110000001111000010111010111111111111100011111111;
    wire [5:0] lut_58_select = {
                             in_data[1143],
                             in_data[2109],
                             in_data[1790],
                             in_data[957],
                             in_data[463],
                             in_data[1697]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [63:0] lut_59_table = 64'b1101111110000001110011010000011111011111000000011100010100000000;
    wire [5:0] lut_59_select = {
                             in_data[655],
                             in_data[704],
                             in_data[746],
                             in_data[1632],
                             in_data[1757],
                             in_data[1113]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [63:0] lut_60_table = 64'b0000000001000000001000000000000011110011111111001011101010111000;
    wire [5:0] lut_60_select = {
                             in_data[785],
                             in_data[703],
                             in_data[1379],
                             in_data[1073],
                             in_data[2111],
                             in_data[1952]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [63:0] lut_61_table = 64'b1111111111110000111111111111111111111111000000001111111101110000;
    wire [5:0] lut_61_select = {
                             in_data[836],
                             in_data[1531],
                             in_data[96],
                             in_data[1232],
                             in_data[136],
                             in_data[544]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [63:0] lut_62_table = 64'b0011000001110000001000001111000011111110111100101110000011110000;
    wire [5:0] lut_62_select = {
                             in_data[2211],
                             in_data[497],
                             in_data[539],
                             in_data[1568],
                             in_data[2268],
                             in_data[1780]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [63:0] lut_63_table = 64'b0000000000000000110111110100111100000000000000101111111111111111;
    wire [5:0] lut_63_select = {
                             in_data[1370],
                             in_data[1373],
                             in_data[102],
                             in_data[792],
                             in_data[1532],
                             in_data[591]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [63:0] lut_64_table = 64'b1111010111000100111111111111110111010100110000001111010111110100;
    wire [5:0] lut_64_select = {
                             in_data[904],
                             in_data[448],
                             in_data[457],
                             in_data[1840],
                             in_data[1694],
                             in_data[985]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [63:0] lut_65_table = 64'b0100001101110001000000001111011100101010000000001111111110110010;
    wire [5:0] lut_65_select = {
                             in_data[1782],
                             in_data[2243],
                             in_data[1740],
                             in_data[1109],
                             in_data[1753],
                             in_data[2174]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [63:0] lut_66_table = 64'b1000100000000000110001000100000011001100000000001111110011111010;
    wire [5:0] lut_66_select = {
                             in_data[1218],
                             in_data[573],
                             in_data[1652],
                             in_data[1380],
                             in_data[568],
                             in_data[2205]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [63:0] lut_67_table = 64'b1101111111011111110111111101111111001111110011001101111101011111;
    wire [5:0] lut_67_select = {
                             in_data[1596],
                             in_data[391],
                             in_data[410],
                             in_data[1789],
                             in_data[1165],
                             in_data[2060]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [63:0] lut_68_table = 64'b1110101011111011110011001100111111111000110010100100110000001100;
    wire [5:0] lut_68_select = {
                             in_data[2252],
                             in_data[1016],
                             in_data[1801],
                             in_data[516],
                             in_data[260],
                             in_data[2195]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [63:0] lut_69_table = 64'b1110111100000100111001000000010011001111000011111110111011001111;
    wire [5:0] lut_69_select = {
                             in_data[911],
                             in_data[709],
                             in_data[441],
                             in_data[2026],
                             in_data[284],
                             in_data[206]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [63:0] lut_70_table = 64'b1111000001010000111111010111000011110000001100001111111111110011;
    wire [5:0] lut_70_select = {
                             in_data[658],
                             in_data[582],
                             in_data[581],
                             in_data[327],
                             in_data[1705],
                             in_data[1417]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [63:0] lut_71_table = 64'b1100111100001111110011110100111100001111000000000000000000000000;
    wire [5:0] lut_71_select = {
                             in_data[1964],
                             in_data[988],
                             in_data[1994],
                             in_data[764],
                             in_data[732],
                             in_data[758]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [63:0] lut_72_table = 64'b0000111000101111000011110010111100001111001011110000011000101011;
    wire [5:0] lut_72_select = {
                             in_data[1489],
                             in_data[1416],
                             in_data[1758],
                             in_data[324],
                             in_data[1664],
                             in_data[86]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [63:0] lut_73_table = 64'b1010101010101010111011101110111011111100111111111111111011111110;
    wire [5:0] lut_73_select = {
                             in_data[82],
                             in_data[1798],
                             in_data[234],
                             in_data[1665],
                             in_data[1912],
                             in_data[776]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [63:0] lut_74_table = 64'b0011111100111111101111111111111111111111001111111110111100001100;
    wire [5:0] lut_74_select = {
                             in_data[1512],
                             in_data[2078],
                             in_data[2282],
                             in_data[317],
                             in_data[1769],
                             in_data[2161]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [63:0] lut_75_table = 64'b1010101011101110111011111111111110101010110010001010101011101111;
    wire [5:0] lut_75_select = {
                             in_data[2155],
                             in_data[440],
                             in_data[1659],
                             in_data[775],
                             in_data[59],
                             in_data[0]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [63:0] lut_76_table = 64'b1101110111011101000000001100110011001100010001000000000001000100;
    wire [5:0] lut_76_select = {
                             in_data[1362],
                             in_data[401],
                             in_data[69],
                             in_data[1990],
                             in_data[639],
                             in_data[406]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [63:0] lut_77_table = 64'b1011101010101010111100101111101111111110101110111111111111111111;
    wire [5:0] lut_77_select = {
                             in_data[1934],
                             in_data[1808],
                             in_data[62],
                             in_data[673],
                             in_data[325],
                             in_data[1106]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [63:0] lut_78_table = 64'b0101000000010000010100000000000011111111011111111101110101000100;
    wire [5:0] lut_78_select = {
                             in_data[823],
                             in_data[2031],
                             in_data[2024],
                             in_data[1354],
                             in_data[405],
                             in_data[794]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [63:0] lut_79_table = 64'b0111000111110111001100110011001101110000111100000000001000000010;
    wire [5:0] lut_79_select = {
                             in_data[1784],
                             in_data[1961],
                             in_data[492],
                             in_data[865],
                             in_data[1468],
                             in_data[1703]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [63:0] lut_80_table = 64'b1101000111010001000000010001010111000100110001001111010101010101;
    wire [5:0] lut_80_select = {
                             in_data[520],
                             in_data[1910],
                             in_data[670],
                             in_data[2086],
                             in_data[773],
                             in_data[387]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [63:0] lut_81_table = 64'b1111011111111101111111111111110100110011101100111111011111111111;
    wire [5:0] lut_81_select = {
                             in_data[2235],
                             in_data[2080],
                             in_data[2004],
                             in_data[390],
                             in_data[2022],
                             in_data[584]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [63:0] lut_82_table = 64'b1011010111110101101000001000000010100101111101010000000000000100;
    wire [5:0] lut_82_select = {
                             in_data[962],
                             in_data[1158],
                             in_data[11],
                             in_data[453],
                             in_data[693],
                             in_data[864]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [63:0] lut_83_table = 64'b1111000011110101111100001111010111110100111101111101000011110000;
    wire [5:0] lut_83_select = {
                             in_data[647],
                             in_data[1361],
                             in_data[1702],
                             in_data[2021],
                             in_data[293],
                             in_data[1484]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [63:0] lut_84_table = 64'b0000000010101100000000001000000010101000111110101010100011111000;
    wire [5:0] lut_84_select = {
                             in_data[1877],
                             in_data[592],
                             in_data[311],
                             in_data[442],
                             in_data[93],
                             in_data[1718]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [63:0] lut_85_table = 64'b1111010011111101111101001101010011111100111111001111010101010000;
    wire [5:0] lut_85_select = {
                             in_data[1328],
                             in_data[1409],
                             in_data[1244],
                             in_data[2180],
                             in_data[900],
                             in_data[1058]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [63:0] lut_86_table = 64'b1111111111111111111011101110111011111011111010111110000011100000;
    wire [5:0] lut_86_select = {
                             in_data[398],
                             in_data[272],
                             in_data[1562],
                             in_data[2263],
                             in_data[1572],
                             in_data[1050]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [63:0] lut_87_table = 64'b1111111101010111111111110100010101010111010001010101011100000000;
    wire [5:0] lut_87_select = {
                             in_data[2007],
                             in_data[2166],
                             in_data[1638],
                             in_data[1344],
                             in_data[371],
                             in_data[37]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [63:0] lut_88_table = 64'b1011000110110001000000001111100010110011000100010000000000010000;
    wire [5:0] lut_88_select = {
                             in_data[1114],
                             in_data[2193],
                             in_data[607],
                             in_data[1076],
                             in_data[2123],
                             in_data[283]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [63:0] lut_89_table = 64'b1111110011010101100000001101010111111100010101010000100001010100;
    wire [5:0] lut_89_select = {
                             in_data[1674],
                             in_data[2226],
                             in_data[837],
                             in_data[945],
                             in_data[1663],
                             in_data[624]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [63:0] lut_90_table = 64'b0000101011011100001010101111101011111111110111001011101011110000;
    wire [5:0] lut_90_select = {
                             in_data[266],
                             in_data[839],
                             in_data[1066],
                             in_data[295],
                             in_data[1097],
                             in_data[1737]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [63:0] lut_91_table = 64'b1100000000000000111110101111111000100000101000001111101011111010;
    wire [5:0] lut_91_select = {
                             in_data[802],
                             in_data[1317],
                             in_data[1064],
                             in_data[1772],
                             in_data[1942],
                             in_data[1429]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [63:0] lut_92_table = 64'b0000100000001010100010101111111100000000000000000000101010001110;
    wire [5:0] lut_92_select = {
                             in_data[2000],
                             in_data[1271],
                             in_data[1829],
                             in_data[2204],
                             in_data[2063],
                             in_data[1637]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [63:0] lut_93_table = 64'b1010000010100000101000001010000011111010111110111110101010100000;
    wire [5:0] lut_93_select = {
                             in_data[1185],
                             in_data[960],
                             in_data[876],
                             in_data[471],
                             in_data[1277],
                             in_data[1907]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [63:0] lut_94_table = 64'b1100110011101100110011001100110011000100110001001100110011111100;
    wire [5:0] lut_94_select = {
                             in_data[1748],
                             in_data[1289],
                             in_data[2295],
                             in_data[143],
                             in_data[616],
                             in_data[1736]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [63:0] lut_95_table = 64'b0000000000100010101111111010111111010000111111111111111111111111;
    wire [5:0] lut_95_select = {
                             in_data[2120],
                             in_data[731],
                             in_data[1499],
                             in_data[1259],
                             in_data[1298],
                             in_data[1085]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [63:0] lut_96_table = 64'b1111101011100000111110100110000011111111111111111111101011111010;
    wire [5:0] lut_96_select = {
                             in_data[1661],
                             in_data[1191],
                             in_data[32],
                             in_data[150],
                             in_data[2034],
                             in_data[1565]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [63:0] lut_97_table = 64'b0010000000000000000011001000110000110010101000000011101111101111;
    wire [5:0] lut_97_select = {
                             in_data[416],
                             in_data[2044],
                             in_data[1336],
                             in_data[495],
                             in_data[762],
                             in_data[828]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [63:0] lut_98_table = 64'b1011101010100010111101110001000010110011001000000111011100010000;
    wire [5:0] lut_98_select = {
                             in_data[362],
                             in_data[614],
                             in_data[1962],
                             in_data[314],
                             in_data[1131],
                             in_data[1832]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [63:0] lut_99_table = 64'b1000100010101111110010001010101000000000101010101000000010101010;
    wire [5:0] lut_99_select = {
                             in_data[2159],
                             in_data[1451],
                             in_data[1810],
                             in_data[838],
                             in_data[156],
                             in_data[75]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [63:0] lut_100_table = 64'b1111111100000011111111110101000100000000000000001111111101011101;
    wire [5:0] lut_100_select = {
                             in_data[74],
                             in_data[2030],
                             in_data[1207],
                             in_data[1590],
                             in_data[1759],
                             in_data[1584]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [63:0] lut_101_table = 64'b1110111111101111100011101010111111101111111111111110111011111111;
    wire [5:0] lut_101_select = {
                             in_data[1929],
                             in_data[103],
                             in_data[698],
                             in_data[135],
                             in_data[2052],
                             in_data[1117]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [63:0] lut_102_table = 64'b0000000001110000001101110111001100000011111100110000001101110011;
    wire [5:0] lut_102_select = {
                             in_data[824],
                             in_data[1447],
                             in_data[641],
                             in_data[1560],
                             in_data[1519],
                             in_data[835]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [63:0] lut_103_table = 64'b1110111110101111101011001010111110001000101011100000000010101010;
    wire [5:0] lut_103_select = {
                             in_data[2227],
                             in_data[1615],
                             in_data[1261],
                             in_data[2220],
                             in_data[800],
                             in_data[885]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [63:0] lut_104_table = 64'b1111111100000111111111110000011100000011000000000111111100000001;
    wire [5:0] lut_104_select = {
                             in_data[235],
                             in_data[2202],
                             in_data[1228],
                             in_data[558],
                             in_data[2125],
                             in_data[1142]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [63:0] lut_105_table = 64'b0000000000000101000001010101010100000000000000000000000000000000;
    wire [5:0] lut_105_select = {
                             in_data[496],
                             in_data[1198],
                             in_data[1792],
                             in_data[553],
                             in_data[127],
                             in_data[194]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [63:0] lut_106_table = 64'b0011000010110010111111111111111100110000001000001111001111111010;
    wire [5:0] lut_106_select = {
                             in_data[515],
                             in_data[1900],
                             in_data[915],
                             in_data[87],
                             in_data[929],
                             in_data[1490]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [63:0] lut_107_table = 64'b0001001100011101000000010000000100111011011111110011001101111111;
    wire [5:0] lut_107_select = {
                             in_data[1860],
                             in_data[1677],
                             in_data[1223],
                             in_data[498],
                             in_data[2113],
                             in_data[240]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [63:0] lut_108_table = 64'b1111101011111010111110111011101011110000101000101111101111111010;
    wire [5:0] lut_108_select = {
                             in_data[569],
                             in_data[716],
                             in_data[2046],
                             in_data[1613],
                             in_data[1184],
                             in_data[1202]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [63:0] lut_109_table = 64'b0111011111111111001100110111011100010000111111110011000101010101;
    wire [5:0] lut_109_select = {
                             in_data[722],
                             in_data[917],
                             in_data[556],
                             in_data[36],
                             in_data[72],
                             in_data[115]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [63:0] lut_110_table = 64'b1111110101110100111111010101000011111111010101001111111100000000;
    wire [5:0] lut_110_select = {
                             in_data[1024],
                             in_data[734],
                             in_data[2106],
                             in_data[955],
                             in_data[438],
                             in_data[273]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [63:0] lut_111_table = 64'b0000001101010101000100010101010100000011000000000010001100000011;
    wire [5:0] lut_111_select = {
                             in_data[1505],
                             in_data[124],
                             in_data[259],
                             in_data[2209],
                             in_data[430],
                             in_data[2057]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [63:0] lut_112_table = 64'b0000000000000000001000100011001100100010010101011010101001110111;
    wire [5:0] lut_112_select = {
                             in_data[2083],
                             in_data[2101],
                             in_data[798],
                             in_data[2239],
                             in_data[1573],
                             in_data[1914]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [63:0] lut_113_table = 64'b1100111100001110100010101000100001011111000111111000101110100010;
    wire [5:0] lut_113_select = {
                             in_data[2029],
                             in_data[1711],
                             in_data[1776],
                             in_data[1850],
                             in_data[157],
                             in_data[80]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [63:0] lut_114_table = 64'b0011111111111100010111111100110000111011000111000011111100001000;
    wire [5:0] lut_114_select = {
                             in_data[2077],
                             in_data[1474],
                             in_data[1141],
                             in_data[1500],
                             in_data[968],
                             in_data[153]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [63:0] lut_115_table = 64'b1110000010111111111100001111011100000000111100111100000011110011;
    wire [5:0] lut_115_select = {
                             in_data[2303],
                             in_data[1744],
                             in_data[1315],
                             in_data[1996],
                             in_data[1537],
                             in_data[1650]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [63:0] lut_116_table = 64'b1111111110001010110011110000000011111101111011101101110011000000;
    wire [5:0] lut_116_select = {
                             in_data[1196],
                             in_data[1092],
                             in_data[1212],
                             in_data[1551],
                             in_data[685],
                             in_data[275]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [63:0] lut_117_table = 64'b0101000011111101010100001111110111110100111111111111000011111100;
    wire [5:0] lut_117_select = {
                             in_data[546],
                             in_data[760],
                             in_data[1025],
                             in_data[799],
                             in_data[594],
                             in_data[1017]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [63:0] lut_118_table = 64'b1010111100000010001010100000001010111111001011111011111100101011;
    wire [5:0] lut_118_select = {
                             in_data[612],
                             in_data[2293],
                             in_data[1817],
                             in_data[1570],
                             in_data[1571],
                             in_data[1793]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [63:0] lut_119_table = 64'b0000111111011111000010010000110100001011010011010000111101011111;
    wire [5:0] lut_119_select = {
                             in_data[645],
                             in_data[1038],
                             in_data[1825],
                             in_data[1339],
                             in_data[285],
                             in_data[2272]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [63:0] lut_120_table = 64'b0101010101001101000000010000100001010101010001010000000000000000;
    wire [5:0] lut_120_select = {
                             in_data[425],
                             in_data[241],
                             in_data[1313],
                             in_data[1217],
                             in_data[1486],
                             in_data[1689]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [63:0] lut_121_table = 64'b0000000000000000100010001000100000001110000000001111111011001000;
    wire [5:0] lut_121_select = {
                             in_data[644],
                             in_data[1267],
                             in_data[38],
                             in_data[843],
                             in_data[2206],
                             in_data[2257]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [63:0] lut_122_table = 64'b1111111101111111011111110000011101111111000001110000011100000111;
    wire [5:0] lut_122_select = {
                             in_data[1641],
                             in_data[643],
                             in_data[264],
                             in_data[1367],
                             in_data[807],
                             in_data[872]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [63:0] lut_123_table = 64'b1010100011111111000000001110111110000000111111110000000010001100;
    wire [5:0] lut_123_select = {
                             in_data[1055],
                             in_data[1986],
                             in_data[1054],
                             in_data[1712],
                             in_data[1540],
                             in_data[708]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [63:0] lut_124_table = 64'b0000111100111010001110110011101000001111000011100011111110111010;
    wire [5:0] lut_124_select = {
                             in_data[1372],
                             in_data[2076],
                             in_data[145],
                             in_data[2027],
                             in_data[477],
                             in_data[354]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [63:0] lut_125_table = 64'b1111111110001111000000000000000011111111101111110010001100000010;
    wire [5:0] lut_125_select = {
                             in_data[1746],
                             in_data[1886],
                             in_data[1049],
                             in_data[998],
                             in_data[1004],
                             in_data[1504]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [63:0] lut_126_table = 64'b1100010011110111000000000101010110000000110101010000000000000000;
    wire [5:0] lut_126_select = {
                             in_data[47],
                             in_data[735],
                             in_data[2146],
                             in_data[1634],
                             in_data[24],
                             in_data[197]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [63:0] lut_127_table = 64'b1000100011001100000000001101111111001111010011010000010011011111;
    wire [5:0] lut_127_select = {
                             in_data[1098],
                             in_data[159],
                             in_data[613],
                             in_data[2012],
                             in_data[855],
                             in_data[1262]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [63:0] lut_128_table = 64'b0000000100000000001000110010001100000011001000110011011100101111;
    wire [5:0] lut_128_select = {
                             in_data[1956],
                             in_data[2278],
                             in_data[525],
                             in_data[631],
                             in_data[1177],
                             in_data[356]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [63:0] lut_129_table = 64'b0101000000001010010101010000000001010010000010100101010100001010;
    wire [5:0] lut_129_select = {
                             in_data[1872],
                             in_data[88],
                             in_data[348],
                             in_data[2126],
                             in_data[2038],
                             in_data[1057]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [63:0] lut_130_table = 64'b0000111100001111001111110000111100001111000011110011111100001111;
    wire [5:0] lut_130_select = {
                             in_data[220],
                             in_data[1645],
                             in_data[1691],
                             in_data[1335],
                             in_data[2185],
                             in_data[766]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [63:0] lut_131_table = 64'b1000111100000000110011110000111010001111000001001100111100000100;
    wire [5:0] lut_131_select = {
                             in_data[2183],
                             in_data[1423],
                             in_data[1545],
                             in_data[931],
                             in_data[1647],
                             in_data[42]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [63:0] lut_132_table = 64'b1011100010111010111110111011101110110000001000101011101100110010;
    wire [5:0] lut_132_select = {
                             in_data[2036],
                             in_data[1670],
                             in_data[1460],
                             in_data[2260],
                             in_data[1378],
                             in_data[1530]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [63:0] lut_133_table = 64'b1100010011110101010011001111110111111101111101110000010000000101;
    wire [5:0] lut_133_select = {
                             in_data[316],
                             in_data[301],
                             in_data[1853],
                             in_data[2276],
                             in_data[1205],
                             in_data[1640]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [63:0] lut_134_table = 64'b0100111011111111110010001100110011001111010111111100110011001100;
    wire [5:0] lut_134_select = {
                             in_data[413],
                             in_data[41],
                             in_data[813],
                             in_data[869],
                             in_data[216],
                             in_data[1461]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [63:0] lut_135_table = 64'b0000000000000000000100000101110100000000000100000001000001010001;
    wire [5:0] lut_135_select = {
                             in_data[626],
                             in_data[1051],
                             in_data[599],
                             in_data[73],
                             in_data[1699],
                             in_data[1148]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [63:0] lut_136_table = 64'b1111111111111111110111001101010011111111000000001101110000000000;
    wire [5:0] lut_136_select = {
                             in_data[1549],
                             in_data[825],
                             in_data[1704],
                             in_data[119],
                             in_data[1709],
                             in_data[1725]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [63:0] lut_137_table = 64'b0000000011111111000000001010101010100000111011100000000011101100;
    wire [5:0] lut_137_select = {
                             in_data[1231],
                             in_data[1760],
                             in_data[826],
                             in_data[1507],
                             in_data[1927],
                             in_data[534]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [63:0] lut_138_table = 64'b1000111011111111100011111111111100001010000000000000101010101110;
    wire [5:0] lut_138_select = {
                             in_data[5],
                             in_data[2059],
                             in_data[2264],
                             in_data[848],
                             in_data[1535],
                             in_data[2068]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [63:0] lut_139_table = 64'b1110011111101111111001110010010011100110111001101110001001100110;
    wire [5:0] lut_139_select = {
                             in_data[1019],
                             in_data[1034],
                             in_data[1954],
                             in_data[1617],
                             in_data[682],
                             in_data[842]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [63:0] lut_140_table = 64'b0000111100001111000111111011111100001111000011110000111110011111;
    wire [5:0] lut_140_select = {
                             in_data[979],
                             in_data[1745],
                             in_data[464],
                             in_data[91],
                             in_data[343],
                             in_data[767]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [63:0] lut_141_table = 64'b0000110100001100010011110000110100000000000000000000110100001000;
    wire [5:0] lut_141_select = {
                             in_data[429],
                             in_data[1115],
                             in_data[474],
                             in_data[597],
                             in_data[550],
                             in_data[1321]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [63:0] lut_142_table = 64'b0101010011001101011101111110111000000000110011110010101010101010;
    wire [5:0] lut_142_select = {
                             in_data[2143],
                             in_data[1435],
                             in_data[2061],
                             in_data[2033],
                             in_data[50],
                             in_data[1681]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [63:0] lut_143_table = 64'b1110100011101000111010001110101011101000111011101110101011101110;
    wire [5:0] lut_143_select = {
                             in_data[681],
                             in_data[1522],
                             in_data[450],
                             in_data[310],
                             in_data[2229],
                             in_data[380]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [63:0] lut_144_table = 64'b0010001000000000111111111111111000110011000000101111111111111111;
    wire [5:0] lut_144_select = {
                             in_data[791],
                             in_data[1696],
                             in_data[1065],
                             in_data[57],
                             in_data[257],
                             in_data[2273]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [63:0] lut_145_table = 64'b0000110000001100111111111110111000001101000011001011111100100010;
    wire [5:0] lut_145_select = {
                             in_data[485],
                             in_data[1386],
                             in_data[137],
                             in_data[784],
                             in_data[454],
                             in_data[331]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [63:0] lut_146_table = 64'b1101100000000000110111011100110111011111110111111101110111011101;
    wire [5:0] lut_146_select = {
                             in_data[2177],
                             in_data[1859],
                             in_data[1951],
                             in_data[2105],
                             in_data[1843],
                             in_data[218]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [63:0] lut_147_table = 64'b0000000000111111000101110011111100000100000111110000010100001111;
    wire [5:0] lut_147_select = {
                             in_data[2224],
                             in_data[1849],
                             in_data[1755],
                             in_data[2279],
                             in_data[595],
                             in_data[1960]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [63:0] lut_148_table = 64'b1011111110111111111110111111111100101011101010100011000010111001;
    wire [5:0] lut_148_select = {
                             in_data[1428],
                             in_data[1015],
                             in_data[951],
                             in_data[1160],
                             in_data[422],
                             in_data[261]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [63:0] lut_149_table = 64'b0000110001001111010101010001000100001100010011110101010101010101;
    wire [5:0] lut_149_select = {
                             in_data[2042],
                             in_data[860],
                             in_data[1786],
                             in_data[1800],
                             in_data[1649],
                             in_data[2085]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [63:0] lut_150_table = 64'b1100110001001100000001010000000001001100110011000100110010001000;
    wire [5:0] lut_150_select = {
                             in_data[1001],
                             in_data[45],
                             in_data[586],
                             in_data[740],
                             in_data[1879],
                             in_data[1145]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [63:0] lut_151_table = 64'b1111110101000100111111011100010011000100110001001100010011000000;
    wire [5:0] lut_151_select = {
                             in_data[65],
                             in_data[801],
                             in_data[1508],
                             in_data[1858],
                             in_data[971],
                             in_data[357]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [63:0] lut_152_table = 64'b0011101000111010000110100011101000001010000010100000101000001110;
    wire [5:0] lut_152_select = {
                             in_data[691],
                             in_data[2280],
                             in_data[1174],
                             in_data[1904],
                             in_data[462],
                             in_data[2259]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [63:0] lut_153_table = 64'b1010100011111011000000001011100010110000101110101010000010110000;
    wire [5:0] lut_153_select = {
                             in_data[176],
                             in_data[672],
                             in_data[1243],
                             in_data[1374],
                             in_data[816],
                             in_data[1511]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [63:0] lut_154_table = 64'b0011111101111111000011111111111100001111011111110000101000111011;
    wire [5:0] lut_154_select = {
                             in_data[227],
                             in_data[26],
                             in_data[48],
                             in_data[744],
                             in_data[547],
                             in_data[1081]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [63:0] lut_155_table = 64'b0000001100000011000100110011001100010011000000110111011101111111;
    wire [5:0] lut_155_select = {
                             in_data[1375],
                             in_data[2006],
                             in_data[2171],
                             in_data[1861],
                             in_data[489],
                             in_data[2066]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [63:0] lut_156_table = 64'b0011000100011111011100010001111111110001000100110001000000010001;
    wire [5:0] lut_156_select = {
                             in_data[1266],
                             in_data[192],
                             in_data[428],
                             in_data[15],
                             in_data[1555],
                             in_data[397]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [63:0] lut_157_table = 64'b0001000000110111000001000001011100001100011111110000110001011111;
    wire [5:0] lut_157_select = {
                             in_data[1846],
                             in_data[1895],
                             in_data[3],
                             in_data[349],
                             in_data[1936],
                             in_data[965]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [63:0] lut_158_table = 64'b0001000001110001000000000111000101001111111111110000000011001111;
    wire [5:0] lut_158_select = {
                             in_data[2090],
                             in_data[1579],
                             in_data[214],
                             in_data[421],
                             in_data[1518],
                             in_data[2160]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [63:0] lut_159_table = 64'b1111111110111111111111111111111100000000000000001111110011111000;
    wire [5:0] lut_159_select = {
                             in_data[878],
                             in_data[207],
                             in_data[1387],
                             in_data[345],
                             in_data[1235],
                             in_data[1981]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [63:0] lut_160_table = 64'b1110111111111111111011110000111110101111101011110010101000001011;
    wire [5:0] lut_160_select = {
                             in_data[1546],
                             in_data[1157],
                             in_data[680],
                             in_data[222],
                             in_data[1329],
                             in_data[1061]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [63:0] lut_161_table = 64'b0001000100000000111100010001000000110001000000001111010100000000;
    wire [5:0] lut_161_select = {
                             in_data[1686],
                             in_data[2158],
                             in_data[251],
                             in_data[654],
                             in_data[1467],
                             in_data[1536]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [63:0] lut_162_table = 64'b1100110011111010110000001000000011011100111111111101010011110001;
    wire [5:0] lut_162_select = {
                             in_data[486],
                             in_data[1881],
                             in_data[262],
                             in_data[519],
                             in_data[1269],
                             in_data[1707]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [63:0] lut_163_table = 64'b1010111000101010101011100010101000101010000000100000101000000010;
    wire [5:0] lut_163_select = {
                             in_data[1195],
                             in_data[25],
                             in_data[867],
                             in_data[1958],
                             in_data[541],
                             in_data[1989]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [63:0] lut_164_table = 64'b0000000000000000111111001100110011001000100010001111110011111110;
    wire [5:0] lut_164_select = {
                             in_data[89],
                             in_data[684],
                             in_data[871],
                             in_data[289],
                             in_data[1525],
                             in_data[2251]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [63:0] lut_165_table = 64'b1111111111011101110011100100111111110101000001010101110100000100;
    wire [5:0] lut_165_select = {
                             in_data[1473],
                             in_data[2092],
                             in_data[19],
                             in_data[1476],
                             in_data[1916],
                             in_data[1974]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [63:0] lut_166_table = 64'b1110111100001110111010100000111000111011000000111111111100110111;
    wire [5:0] lut_166_select = {
                             in_data[1247],
                             in_data[282],
                             in_data[2266],
                             in_data[947],
                             in_data[1820],
                             in_data[1175]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [63:0] lut_167_table = 64'b1101010001010001110011100100011101010010010100110100101000100010;
    wire [5:0] lut_167_select = {
                             in_data[1660],
                             in_data[892],
                             in_data[1639],
                             in_data[563],
                             in_data[532],
                             in_data[2117]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [63:0] lut_168_table = 64'b1111111110101010111011011110000011111111101011111100111110101010;
    wire [5:0] lut_168_select = {
                             in_data[2133],
                             in_data[1411],
                             in_data[1011],
                             in_data[1006],
                             in_data[1236],
                             in_data[1804]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [63:0] lut_169_table = 64'b0000000010000000000000000000000010101110111011111000111011101111;
    wire [5:0] lut_169_select = {
                             in_data[237],
                             in_data[1785],
                             in_data[1287],
                             in_data[1128],
                             in_data[85],
                             in_data[1919]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [63:0] lut_170_table = 64'b1000101011101111000000101000111111101011111111111011101111111111;
    wire [5:0] lut_170_select = {
                             in_data[2148],
                             in_data[2228],
                             in_data[404],
                             in_data[1090],
                             in_data[2269],
                             in_data[1099]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [63:0] lut_171_table = 64'b0011011100000000010101011101110101110111000001001111111111011101;
    wire [5:0] lut_171_select = {
                             in_data[139],
                             in_data[279],
                             in_data[1478],
                             in_data[605],
                             in_data[1342],
                             in_data[2201]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [63:0] lut_172_table = 64'b1101110011111111110001001111110000000000110001000100000011110000;
    wire [5:0] lut_172_select = {
                             in_data[452],
                             in_data[1601],
                             in_data[1643],
                             in_data[1324],
                             in_data[2015],
                             in_data[1233]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [63:0] lut_173_table = 64'b0111001111110111011101111111011101110010011100110111001101110000;
    wire [5:0] lut_173_select = {
                             in_data[389],
                             in_data[1028],
                             in_data[1048],
                             in_data[1014],
                             in_data[449],
                             in_data[974]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [63:0] lut_174_table = 64'b1111111111001111110011101100110011111111110001001000100000000000;
    wire [5:0] lut_174_select = {
                             in_data[656],
                             in_data[724],
                             in_data[300],
                             in_data[1687],
                             in_data[1657],
                             in_data[662]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [63:0] lut_175_table = 64'b1000110111100100000001011100010010001111111111111010111111111111;
    wire [5:0] lut_175_select = {
                             in_data[712],
                             in_data[1220],
                             in_data[690],
                             in_data[2169],
                             in_data[215],
                             in_data[1470]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [63:0] lut_176_table = 64'b1111011111110011111101111111001110100000101100111111000011110010;
    wire [5:0] lut_176_select = {
                             in_data[1834],
                             in_data[1359],
                             in_data[996],
                             in_data[270],
                             in_data[346],
                             in_data[1039]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [63:0] lut_177_table = 64'b0010001000100010001100101011001010111011101010101011101110111011;
    wire [5:0] lut_177_select = {
                             in_data[606],
                             in_data[1706],
                             in_data[1723],
                             in_data[2179],
                             in_data[743],
                             in_data[1306]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [63:0] lut_178_table = 64'b0010111110101111001000111011111100000101000111110000000000000001;
    wire [5:0] lut_178_select = {
                             in_data[665],
                             in_data[2035],
                             in_data[632],
                             in_data[1625],
                             in_data[2091],
                             in_data[1865]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [63:0] lut_179_table = 64'b0000111100010101000011110000110100000111000001010000111100000100;
    wire [5:0] lut_179_select = {
                             in_data[294],
                             in_data[1612],
                             in_data[804],
                             in_data[1675],
                             in_data[2246],
                             in_data[529]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [63:0] lut_180_table = 64'b0000000000000000010101010000010111111111000001011111111100000101;
    wire [5:0] lut_180_select = {
                             in_data[1575],
                             in_data[609],
                             in_data[1813],
                             in_data[1042],
                             in_data[195],
                             in_data[1010]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [63:0] lut_181_table = 64'b0000000000001100000011000000111100000100000011011000111100111111;
    wire [5:0] lut_181_select = {
                             in_data[376],
                             in_data[1360],
                             in_data[1187],
                             in_data[946],
                             in_data[1035],
                             in_data[1585]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [63:0] lut_182_table = 64'b1111111100001000111111110000100011001100000000001101111100000101;
    wire [5:0] lut_182_select = {
                             in_data[1925],
                             in_data[870],
                             in_data[2050],
                             in_data[1690],
                             in_data[437],
                             in_data[27]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [63:0] lut_183_table = 64'b1111001011111000111110111111101111110001110100001111001111111011;
    wire [5:0] lut_183_select = {
                             in_data[2054],
                             in_data[2055],
                             in_data[71],
                             in_data[2164],
                             in_data[1902],
                             in_data[263]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [63:0] lut_184_table = 64'b1111010011000000111100000000000011111110111010101111111011101111;
    wire [5:0] lut_184_select = {
                             in_data[1984],
                             in_data[493],
                             in_data[1116],
                             in_data[1393],
                             in_data[718],
                             in_data[1869]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [63:0] lut_185_table = 64'b0000010100000101000010000000100001000101010011111010111010101110;
    wire [5:0] lut_185_select = {
                             in_data[483],
                             in_data[1291],
                             in_data[372],
                             in_data[1107],
                             in_data[883],
                             in_data[1855]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [63:0] lut_186_table = 64'b0011001100100010001000110010001100000000001000001011101100101011;
    wire [5:0] lut_186_select = {
                             in_data[728],
                             in_data[287],
                             in_data[1304],
                             in_data[304],
                             in_data[1343],
                             in_data[1947]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [63:0] lut_187_table = 64'b0001011100000001000101110001011100011111000101011111111111111101;
    wire [5:0] lut_187_select = {
                             in_data[487],
                             in_data[714],
                             in_data[1826],
                             in_data[1334],
                             in_data[899],
                             in_data[610]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [63:0] lut_188_table = 64'b0000101000001010000010000000000011101111111111111111111111001010;
    wire [5:0] lut_188_select = {
                             in_data[1465],
                             in_data[1087],
                             in_data[219],
                             in_data[964],
                             in_data[922],
                             in_data[1618]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [63:0] lut_189_table = 64'b0000000011111111000010001111111110101000111111110010000011111111;
    wire [5:0] lut_189_select = {
                             in_data[1176],
                             in_data[747],
                             in_data[1462],
                             in_data[1154],
                             in_data[180],
                             in_data[981]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [63:0] lut_190_table = 64'b0100010000000000011101000000000011011100000001001111110100000100;
    wire [5:0] lut_190_select = {
                             in_data[17],
                             in_data[2289],
                             in_data[1250],
                             in_data[1581],
                             in_data[2132],
                             in_data[1965]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [63:0] lut_191_table = 64'b1101110111000100111100001101000011001111110010011111111111000001;
    wire [5:0] lut_191_select = {
                             in_data[2254],
                             in_data[1316],
                             in_data[2151],
                             in_data[1404],
                             in_data[1610],
                             in_data[2043]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [63:0] lut_192_table = 64'b1011101111011100000000001101110000000000100000001101000011111100;
    wire [5:0] lut_192_select = {
                             in_data[66],
                             in_data[1418],
                             in_data[897],
                             in_data[1837],
                             in_data[2299],
                             in_data[455]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [63:0] lut_193_table = 64'b1111011110100011011100010001000011111111011111111111011100000001;
    wire [5:0] lut_193_select = {
                             in_data[1970],
                             in_data[199],
                             in_data[577],
                             in_data[719],
                             in_data[1903],
                             in_data[2124]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [63:0] lut_194_table = 64'b1111111111111111100000000000000011111110111101110000101000000000;
    wire [5:0] lut_194_select = {
                             in_data[323],
                             in_data[1897],
                             in_data[1285],
                             in_data[687],
                             in_data[1458],
                             in_data[35]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [63:0] lut_195_table = 64'b1111100011111010111111111111111100000000000000000101010001010001;
    wire [5:0] lut_195_select = {
                             in_data[1299],
                             in_data[2023],
                             in_data[1972],
                             in_data[461],
                             in_data[642],
                             in_data[621]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [63:0] lut_196_table = 64'b0001010111010000000000110101000000010111010101010001001101010001;
    wire [5:0] lut_196_select = {
                             in_data[1211],
                             in_data[2285],
                             in_data[858],
                             in_data[1620],
                             in_data[407],
                             in_data[1475]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [63:0] lut_197_table = 64'b1001000011010001000100000001000111011101111111110101000111011101;
    wire [5:0] lut_197_select = {
                             in_data[2065],
                             in_data[1063],
                             in_data[1410],
                             in_data[1003],
                             in_data[303],
                             in_data[394]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [63:0] lut_198_table = 64'b0100010001001100000001000100010000000000000000000000000000000000;
    wire [5:0] lut_198_select = {
                             in_data[433],
                             in_data[92],
                             in_data[347],
                             in_data[1741],
                             in_data[874],
                             in_data[575]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [63:0] lut_199_table = 64'b0010000000000000101100110011001010110010101100000010000000100000;
    wire [5:0] lut_199_select = {
                             in_data[1279],
                             in_data[1353],
                             in_data[183],
                             in_data[1406],
                             in_data[753],
                             in_data[144]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [63:0] lut_200_table = 64'b0000000000100010000000000010001110101011101110100010001000101010;
    wire [5:0] lut_200_select = {
                             in_data[2016],
                             in_data[588],
                             in_data[1056],
                             in_data[202],
                             in_data[276],
                             in_data[1371]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [63:0] lut_201_table = 64'b0010101100000010101011110000001110100011000000111010101100000011;
    wire [5:0] lut_201_select = {
                             in_data[1290],
                             in_data[1095],
                             in_data[1403],
                             in_data[95],
                             in_data[1944],
                             in_data[821]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [63:0] lut_202_table = 64'b1000111011001100000010100000111111111111111111001111111111111111;
    wire [5:0] lut_202_select = {
                             in_data[205],
                             in_data[2262],
                             in_data[1273],
                             in_data[2144],
                             in_data[2095],
                             in_data[30]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [63:0] lut_203_table = 64'b1111111111001111110011110000110011111111111111111100111111001100;
    wire [5:0] lut_203_select = {
                             in_data[2294],
                             in_data[196],
                             in_data[862],
                             in_data[1662],
                             in_data[189],
                             in_data[1036]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [63:0] lut_204_table = 64'b1010101010101010100010001010100010101000101110101000000010111000;
    wire [5:0] lut_204_select = {
                             in_data[1144],
                             in_data[411],
                             in_data[439],
                             in_data[1513],
                             in_data[107],
                             in_data[1523]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [63:0] lut_205_table = 64'b0011001100110011011100000011000000110000001100001111000011110000;
    wire [5:0] lut_205_select = {
                             in_data[1909],
                             in_data[1483],
                             in_data[1255],
                             in_data[247],
                             in_data[1594],
                             in_data[1949]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [63:0] lut_206_table = 64'b0101111101001101010111110100010111110011001100110001000100010001;
    wire [5:0] lut_206_select = {
                             in_data[806],
                             in_data[651],
                             in_data[786],
                             in_data[1121],
                             in_data[1162],
                             in_data[694]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [63:0] lut_207_table = 64'b1101111011111111000000001000101011111100111111110100000011000010;
    wire [5:0] lut_207_select = {
                             in_data[1307],
                             in_data[379],
                             in_data[1469],
                             in_data[181],
                             in_data[1169],
                             in_data[1534]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [63:0] lut_208_table = 64'b1111111111110111111111111111111111111111000000011111111100000000;
    wire [5:0] lut_208_select = {
                             in_data[1224],
                             in_data[938],
                             in_data[788],
                             in_data[1700],
                             in_data[1922],
                             in_data[1816]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [63:0] lut_209_table = 64'b0000000000000000000000000000110000000000000000001000100011001100;
    wire [5:0] lut_209_select = {
                             in_data[997],
                             in_data[236],
                             in_data[1828],
                             in_data[182],
                             in_data[1779],
                             in_data[2198]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [63:0] lut_210_table = 64'b0000101000001100100010101110111010101110110011101110111011111111;
    wire [5:0] lut_210_select = {
                             in_data[1626],
                             in_data[507],
                             in_data[174],
                             in_data[1971],
                             in_data[120],
                             in_data[420]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [63:0] lut_211_table = 64'b1111001111110010101100111111001010110000111100000000000010100000;
    wire [5:0] lut_211_select = {
                             in_data[61],
                             in_data[1874],
                             in_data[2241],
                             in_data[926],
                             in_data[866],
                             in_data[741]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [63:0] lut_212_table = 64'b0001000011111100011111111111111100000000000000000000001000110010;
    wire [5:0] lut_212_select = {
                             in_data[226],
                             in_data[1501],
                             in_data[761],
                             in_data[1413],
                             in_data[840],
                             in_data[1348]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [63:0] lut_213_table = 64'b0000000100000111000000110001111100000000000000000000000001011111;
    wire [5:0] lut_213_select = {
                             in_data[1407],
                             in_data[528],
                             in_data[187],
                             in_data[1482],
                             in_data[79],
                             in_data[1292]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [63:0] lut_214_table = 64'b1111111100101111111011111110111100001111000001110000001100000011;
    wire [5:0] lut_214_select = {
                             in_data[1997],
                             in_data[459],
                             in_data[557],
                             in_data[1926],
                             in_data[1147],
                             in_data[552]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [63:0] lut_215_table = 64'b0000100000101011000011110011111100000000001010110000000000100011;
    wire [5:0] lut_215_select = {
                             in_data[1319],
                             in_data[2223],
                             in_data[110],
                             in_data[31],
                             in_data[841],
                             in_data[720]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [63:0] lut_216_table = 64'b0011111100000111111111110001111100000000000000000000001100000000;
    wire [5:0] lut_216_select = {
                             in_data[426],
                             in_data[435],
                             in_data[434],
                             in_data[1498],
                             in_data[1448],
                             in_data[1264]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [63:0] lut_217_table = 64'b0000110011001101000111111111111100000000010000000001001111010001;
    wire [5:0] lut_217_select = {
                             in_data[1268],
                             in_data[664],
                             in_data[939],
                             in_data[1083],
                             in_data[1905],
                             in_data[1040]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [63:0] lut_218_table = 64'b0011001111111111000000001111011100110011111100110111011111111111;
    wire [5:0] lut_218_select = {
                             in_data[1186],
                             in_data[1401],
                             in_data[2238],
                             in_data[928],
                             in_data[277],
                             in_data[1449]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [63:0] lut_219_table = 64'b1110111111001100101000000000000010101111111111111010001100110111;
    wire [5:0] lut_219_select = {
                             in_data[1341],
                             in_data[1368],
                             in_data[1633],
                             in_data[567],
                             in_data[258],
                             in_data[1093]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [63:0] lut_220_table = 64'b1110100000100000101111110000000010100000000000000000000100000000;
    wire [5:0] lut_220_select = {
                             in_data[1515],
                             in_data[1685],
                             in_data[1112],
                             in_data[1667],
                             in_data[305],
                             in_data[908]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [63:0] lut_221_table = 64'b0000111101010111010011110000010110101111111111111010111100000111;
    wire [5:0] lut_221_select = {
                             in_data[1976],
                             in_data[44],
                             in_data[653],
                             in_data[1033],
                             in_data[2037],
                             in_data[1312]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [63:0] lut_222_table = 64'b0101010001010100010000000100010011110100111111110000000000000100;
    wire [5:0] lut_222_select = {
                             in_data[697],
                             in_data[378],
                             in_data[1722],
                             in_data[10],
                             in_data[1778],
                             in_data[2097]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [63:0] lut_223_table = 64'b1111111111001100010000000000000011111111110011110100000000000000;
    wire [5:0] lut_223_select = {
                             in_data[1137],
                             in_data[100],
                             in_data[778],
                             in_data[1836],
                             in_data[700],
                             in_data[1756]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [63:0] lut_224_table = 64'b1101111101000100110111110100110011111111000000000001001000000000;
    wire [5:0] lut_224_select = {
                             in_data[23],
                             in_data[2162],
                             in_data[2283],
                             in_data[315],
                             in_data[1108],
                             in_data[1933]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [63:0] lut_225_table = 64'b1111101110110001111110111111101110111011000000001010101010000010;
    wire [5:0] lut_225_select = {
                             in_data[1787],
                             in_data[369],
                             in_data[1521],
                             in_data[1838],
                             in_data[2131],
                             in_data[1636]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [63:0] lut_226_table = 64'b1111110111111101010101000101010100000100110001000000000000000000;
    wire [5:0] lut_226_select = {
                             in_data[733],
                             in_data[388],
                             in_data[1419],
                             in_data[2003],
                             in_data[2222],
                             in_data[1932]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [63:0] lut_227_table = 64'b0101010101000101010001000100010000000010000000100000001000000000;
    wire [5:0] lut_227_select = {
                             in_data[1995],
                             in_data[1946],
                             in_data[559],
                             in_data[1159],
                             in_data[668],
                             in_data[1122]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [63:0] lut_228_table = 64'b0000000000000010001110110010101111000000000000001111111110001110;
    wire [5:0] lut_228_select = {
                             in_data[2119],
                             in_data[2056],
                             in_data[831],
                             in_data[1783],
                             in_data[328],
                             in_data[1999]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [63:0] lut_229_table = 64'b1111011111110111101111111111111100110000011100001011101111111011;
    wire [5:0] lut_229_select = {
                             in_data[1721],
                             in_data[1735],
                             in_data[1364],
                             in_data[383],
                             in_data[446],
                             in_data[99]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [63:0] lut_230_table = 64'b0011000000001100000100000000110000110000000000000011000111111111;
    wire [5:0] lut_230_select = {
                             in_data[1622],
                             in_data[585],
                             in_data[1172],
                             in_data[1078],
                             in_data[1192],
                             in_data[1630]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [63:0] lut_231_table = 64'b0001110100000000010001010000000001011101000001000101010101000100;
    wire [5:0] lut_231_select = {
                             in_data[1682],
                             in_data[1384],
                             in_data[1111],
                             in_data[1992],
                             in_data[1427],
                             in_data[1164]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [63:0] lut_232_table = 64'b1111111010101010111011101010101011101110100010101100111000001110;
    wire [5:0] lut_232_select = {
                             in_data[1219],
                             in_data[1982],
                             in_data[1240],
                             in_data[1213],
                             in_data[1893],
                             in_data[2094]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [63:0] lut_233_table = 64'b0100110101001100010011010000010101001101010011000000010100000101;
    wire [5:0] lut_233_select = {
                             in_data[578],
                             in_data[817],
                             in_data[238],
                             in_data[949],
                             in_data[2053],
                             in_data[1730]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [63:0] lut_234_table = 64'b1101000011010000111100111111000111111000110000001011001111110000;
    wire [5:0] lut_234_select = {
                             in_data[2121],
                             in_data[1953],
                             in_data[832],
                             in_data[1318],
                             in_data[1310],
                             in_data[342]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [63:0] lut_235_table = 64'b0001000000000100000100000001110101010101000011010001000100011101;
    wire [5:0] lut_235_select = {
                             in_data[1577],
                             in_data[1623],
                             in_data[1425],
                             in_data[661],
                             in_data[233],
                             in_data[795]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [63:0] lut_236_table = 64'b1111000011111110111111111111111111100000111100000000000011000000;
    wire [5:0] lut_236_select = {
                             in_data[1864],
                             in_data[1280],
                             in_data[2009],
                             in_data[1492],
                             in_data[280],
                             in_data[975]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [63:0] lut_237_table = 64'b1111110011111101111000001111110011110000111100001111000011110000;
    wire [5:0] lut_237_select = {
                             in_data[1628],
                             in_data[402],
                             in_data[1917],
                             in_data[1203],
                             in_data[877],
                             in_data[686]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [63:0] lut_238_table = 64'b1011001111110111111111111111111100010001011101011011011111111111;
    wire [5:0] lut_238_select = {
                             in_data[1376],
                             in_data[506],
                             in_data[777],
                             in_data[269],
                             in_data[417],
                             in_data[688]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [63:0] lut_239_table = 64'b1111001111110001000000000100000000111111011101110000000000110000;
    wire [5:0] lut_239_select = {
                             in_data[961],
                             in_data[1276],
                             in_data[2140],
                             in_data[1818],
                             in_data[1062],
                             in_data[1493]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [63:0] lut_240_table = 64'b1111101110110010111110101010001010111111000010111011111100001111;
    wire [5:0] lut_240_select = {
                             in_data[1037],
                             in_data[671],
                             in_data[675],
                             in_data[308],
                             in_data[1104],
                             in_data[1765]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [63:0] lut_241_table = 64'b1111011010100010111111101110101000000000101000101000000010101000;
    wire [5:0] lut_241_select = {
                             in_data[1340],
                             in_data[1302],
                             in_data[699],
                             in_data[1574],
                             in_data[1363],
                             in_data[1727]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [63:0] lut_242_table = 64'b1111000000000000111111110000000000000000000000001111111100000000;
    wire [5:0] lut_242_select = {
                             in_data[501],
                             in_data[2087],
                             in_data[781],
                             in_data[706],
                             in_data[1807],
                             in_data[1018]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [63:0] lut_243_table = 64'b1111111100110001111111111111001111110011001100011111111111111011;
    wire [5:0] lut_243_select = {
                             in_data[2082],
                             in_data[1848],
                             in_data[875],
                             in_data[55],
                             in_data[1464],
                             in_data[1139]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [63:0] lut_244_table = 64'b1101110011110101000001000101000011011100111111001100000011010000;
    wire [5:0] lut_244_select = {
                             in_data[1876],
                             in_data[1181],
                             in_data[707],
                             in_data[943],
                             in_data[510],
                             in_data[108]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [63:0] lut_245_table = 64'b1111111111111110000000001111101011111111110111100000100011101010;
    wire [5:0] lut_245_select = {
                             in_data[1602],
                             in_data[1119],
                             in_data[1125],
                             in_data[2073],
                             in_data[2208],
                             in_data[2093]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [63:0] lut_246_table = 64'b0010000000100011000000000000000011111010111011101110100010001000;
    wire [5:0] lut_246_select = {
                             in_data[14],
                             in_data[1242],
                             in_data[2167],
                             in_data[2156],
                             in_data[844],
                             in_data[1957]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [63:0] lut_247_table = 64'b1111111011101010111010101110101011101110101000001010101010100010;
    wire [5:0] lut_247_select = {
                             in_data[1320],
                             in_data[1433],
                             in_data[2290],
                             in_data[1126],
                             in_data[1241],
                             in_data[990]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [63:0] lut_248_table = 64'b0100010111111111010001010101010101010101111111110000010100110111;
    wire [5:0] lut_248_select = {
                             in_data[2072],
                             in_data[1541],
                             in_data[1102],
                             in_data[1136],
                             in_data[2051],
                             in_data[20]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [63:0] lut_249_table = 64'b0010000011110010001000101011001000000000111111110010001011111011;
    wire [5:0] lut_249_select = {
                             in_data[986],
                             in_data[1424],
                             in_data[2267],
                             in_data[910],
                             in_data[488],
                             in_data[51]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [63:0] lut_250_table = 64'b1111000100000000111101110101000101110111000000111101111101000101;
    wire [5:0] lut_250_select = {
                             in_data[1680],
                             in_data[2196],
                             in_data[1132],
                             in_data[1253],
                             in_data[1524],
                             in_data[230]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [63:0] lut_251_table = 64'b0101010101010101000000010100010001010001011101010011000101110101;
    wire [5:0] lut_251_select = {
                             in_data[2118],
                             in_data[576],
                             in_data[166],
                             in_data[1281],
                             in_data[1286],
                             in_data[1284]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [63:0] lut_252_table = 64'b1011111100100011111111100010000010111111001010111010100000000000;
    wire [5:0] lut_252_select = {
                             in_data[1405],
                             in_data[1452],
                             in_data[1338],
                             in_data[2271],
                             in_data[2069],
                             in_data[1889]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [63:0] lut_253_table = 64'b1111111111111111101011110000000000001111000011110000000000000000;
    wire [5:0] lut_253_select = {
                             in_data[1357],
                             in_data[880],
                             in_data[244],
                             in_data[1194],
                             in_data[1988],
                             in_data[705]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [63:0] lut_254_table = 64'b1111001111110011111100111111101100110010000100100011000010110010;
    wire [5:0] lut_254_select = {
                             in_data[958],
                             in_data[1672],
                             in_data[982],
                             in_data[2013],
                             in_data[382],
                             in_data[363]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [63:0] lut_255_table = 64'b1011001000100000111100110000000011110011111100011111111111110011;
    wire [5:0] lut_255_select = {
                             in_data[1210],
                             in_data[168],
                             in_data[560],
                             in_data[1683],
                             in_data[290],
                             in_data[1693]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [63:0] lut_256_table = 64'b0000001110100011001000110011001110101111101011111011111110111111;
    wire [5:0] lut_256_select = {
                             in_data[879],
                             in_data[1987],
                             in_data[1924],
                             in_data[1079],
                             in_data[1450],
                             in_data[414]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [63:0] lut_257_table = 64'b1111000011110000010011011101110111011101111110010101110111111111;
    wire [5:0] lut_257_select = {
                             in_data[846],
                             in_data[2141],
                             in_data[470],
                             in_data[1966],
                             in_data[696],
                             in_data[28]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [63:0] lut_258_table = 64'b1100000000000000000000000000000011111111111010001110110010000000;
    wire [5:0] lut_258_select = {
                             in_data[444],
                             in_data[1878],
                             in_data[2005],
                             in_data[1593],
                             in_data[562],
                             in_data[1152]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [63:0] lut_259_table = 64'b1111111111011111110011110100010110101111101011111000111100001110;
    wire [5:0] lut_259_select = {
                             in_data[123],
                             in_data[738],
                             in_data[1395],
                             in_data[542],
                             in_data[1377],
                             in_data[211]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [63:0] lut_260_table = 64'b0000000100100011000000010010001000000001000101110001000100000001;
    wire [5:0] lut_260_select = {
                             in_data[321],
                             in_data[128],
                             in_data[113],
                             in_data[977],
                             in_data[2084],
                             in_data[1930]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [63:0] lut_261_table = 64'b0000010111111111011111111111111100000111111111110011011111111111;
    wire [5:0] lut_261_select = {
                             in_data[177],
                             in_data[274],
                             in_data[1812],
                             in_data[360],
                             in_data[1294],
                             in_data[424]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [63:0] lut_262_table = 64'b1100110100000000110111110000000011111111010000001111111111110100;
    wire [5:0] lut_262_select = {
                             in_data[1000],
                             in_data[959],
                             in_data[2178],
                             in_data[1631],
                             in_data[1796],
                             in_data[1854]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [63:0] lut_263_table = 64'b1110111111101111011011111110111011001110111011110100110011001100;
    wire [5:0] lut_263_select = {
                             in_data[890],
                             in_data[1044],
                             in_data[140],
                             in_data[148],
                             in_data[1833],
                             in_data[948]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [63:0] lut_264_table = 64'b0010001000001000001000101010000010111010111110101010101011111010;
    wire [5:0] lut_264_select = {
                             in_data[70],
                             in_data[2291],
                             in_data[873],
                             in_data[1870],
                             in_data[491],
                             in_data[1609]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [63:0] lut_265_table = 64'b0111000111110001111110100010001001110000001000001010001000000000;
    wire [5:0] lut_265_select = {
                             in_data[1305],
                             in_data[245],
                             in_data[58],
                             in_data[1075],
                             in_data[278],
                             in_data[1337]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [63:0] lut_266_table = 64'b1100111101001101111111111101111101000100010001001100110011011111;
    wire [5:0] lut_266_select = {
                             in_data[2210],
                             in_data[1496],
                             in_data[1797],
                             in_data[1651],
                             in_data[1863],
                             in_data[891]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [63:0] lut_267_table = 64'b0111000101110101011100000111010000110011011101110001000001110101;
    wire [5:0] lut_267_select = {
                             in_data[352],
                             in_data[271],
                             in_data[351],
                             in_data[1238],
                             in_data[663],
                             in_data[1155]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [63:0] lut_268_table = 64'b1010101010101010101011110000000011101111101000101111111111101111;
    wire [5:0] lut_268_select = {
                             in_data[2275],
                             in_data[1606],
                             in_data[1752],
                             in_data[1383],
                             in_data[1150],
                             in_data[847]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [63:0] lut_269_table = 64'b0000010000000101001001010010010111110111111101110010010100100101;
    wire [5:0] lut_269_select = {
                             in_data[1047],
                             in_data[782],
                             in_data[630],
                             in_data[1008],
                             in_data[618],
                             in_data[1303]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [63:0] lut_270_table = 64'b0000011101110111000000000011000100100000101100110010001010110011;
    wire [5:0] lut_270_select = {
                             in_data[1679],
                             in_data[1739],
                             in_data[1067],
                             in_data[611],
                             in_data[2019],
                             in_data[736]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [63:0] lut_271_table = 64'b0000111100001010001010100000000000001111000011011111110000000000;
    wire [5:0] lut_271_select = {
                             in_data[1552],
                             in_data[1561],
                             in_data[2115],
                             in_data[533],
                             in_data[1365],
                             in_data[1781]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [63:0] lut_272_table = 64'b0111011101011111010101010000010101110111000001010101010100000001;
    wire [5:0] lut_272_select = {
                             in_data[810],
                             in_data[1839],
                             in_data[12],
                             in_data[1347],
                             in_data[231],
                             in_data[1767]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [63:0] lut_273_table = 64'b1111010111011101111101011111010111010101110111011111010111110101;
    wire [5:0] lut_273_select = {
                             in_data[633],
                             in_data[2028],
                             in_data[1012],
                             in_data[118],
                             in_data[1928],
                             in_data[1884]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [63:0] lut_274_table = 64'b0000101100000001111111110001011111111111111111111111111111111111;
    wire [5:0] lut_274_select = {
                             in_data[2129],
                             in_data[2089],
                             in_data[396],
                             in_data[1802],
                             in_data[748],
                             in_data[679]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [63:0] lut_275_table = 64'b0000000000001111000000000000010000001111111011110011110100101111;
    wire [5:0] lut_275_select = {
                             in_data[1480],
                             in_data[2236],
                             in_data[953],
                             in_data[1799],
                             in_data[126],
                             in_data[1091]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [63:0] lut_276_table = 64'b0111010100110000000111110001000001111101001100000110111000001010;
    wire [5:0] lut_276_select = {
                             in_data[1506],
                             in_data[1819],
                             in_data[256],
                             in_data[940],
                             in_data[1],
                             in_data[622]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [63:0] lut_277_table = 64'b0110101111111111000000001110101011011101110011000100110011000000;
    wire [5:0] lut_277_select = {
                             in_data[936],
                             in_data[1455],
                             in_data[105],
                             in_data[2300],
                             in_data[2215],
                             in_data[1844]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [63:0] lut_278_table = 64'b1101010001110100111100001111000011011101001101001111110011111100;
    wire [5:0] lut_278_select = {
                             in_data[1939],
                             in_data[989],
                             in_data[850],
                             in_data[727],
                             in_data[1171],
                             in_data[34]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [63:0] lut_279_table = 64'b0001000011111111000000000000000011111111111111110000101100001010;
    wire [5:0] lut_279_select = {
                             in_data[1221],
                             in_data[505],
                             in_data[768],
                             in_data[1811],
                             in_data[1788],
                             in_data[1005]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [63:0] lut_280_table = 64'b0011001100101011001100110010001100100011000000100010001010100010;
    wire [5:0] lut_280_select = {
                             in_data[755],
                             in_data[353],
                             in_data[1270],
                             in_data[2253],
                             in_data[545],
                             in_data[1434]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [63:0] lut_281_table = 64'b1111001011110010111100101111001011111111111111111111111011111111;
    wire [5:0] lut_281_select = {
                             in_data[659],
                             in_data[1600],
                             in_data[9],
                             in_data[540],
                             in_data[1072],
                             in_data[1724]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [63:0] lut_282_table = 64'b1000111111101111100011001010111110001101101111111011111110111011;
    wire [5:0] lut_282_select = {
                             in_data[1906],
                             in_data[2041],
                             in_data[1118],
                             in_data[1624],
                             in_data[175],
                             in_data[1086]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [63:0] lut_283_table = 64'b1100010001001101110111110100111111110100010100011111010101110111;
    wire [5:0] lut_283_select = {
                             in_data[2207],
                             in_data[178],
                             in_data[593],
                             in_data[395],
                             in_data[500],
                             in_data[1325]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [63:0] lut_284_table = 64'b0001000111010001010000010100000100100011111101011100010111000101;
    wire [5:0] lut_284_select = {
                             in_data[1105],
                             in_data[935],
                             in_data[2079],
                             in_data[2265],
                             in_data[1642],
                             in_data[1188]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [63:0] lut_285_table = 64'b0101110100101011010111110111101100000000000000100001000100000010;
    wire [5:0] lut_285_select = {
                             in_data[1274],
                             in_data[1190],
                             in_data[827],
                             in_data[1237],
                             in_data[881],
                             in_data[375]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [63:0] lut_286_table = 64'b1100000001000000111111001100100011010100010000001111111111001000;
    wire [5:0] lut_286_select = {
                             in_data[933],
                             in_data[590],
                             in_data[2281],
                             in_data[518],
                             in_data[494],
                             in_data[1225]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [63:0] lut_287_table = 64'b0011001110110010001000010010000011110011111100101011000010100000;
    wire [5:0] lut_287_select = {
                             in_data[912],
                             in_data[629],
                             in_data[445],
                             in_data[403],
                             in_data[674],
                             in_data[16]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [63:0] lut_288_table = 64'b1111110000001000111111010000000011111111110011001111110111011100;
    wire [5:0] lut_288_select = {
                             in_data[657],
                             in_data[78],
                             in_data[1582],
                             in_data[1856],
                             in_data[466],
                             in_data[1847]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [63:0] lut_289_table = 64'b0000111101001111000011110000111100001101000011010000111100001111;
    wire [5:0] lut_289_select = {
                             in_data[619],
                             in_data[138],
                             in_data[1134],
                             in_data[2128],
                             in_data[1768],
                             in_data[1227]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [63:0] lut_290_table = 64'b0010101100100010000010110010001011111010111100000010001011110000;
    wire [5:0] lut_290_select = {
                             in_data[104],
                             in_data[1963],
                             in_data[1991],
                             in_data[1481],
                             in_data[1899],
                             in_data[21]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [63:0] lut_291_table = 64'b0000000000001010000010001011101100000000000010100000001110111011;
    wire [5:0] lut_291_select = {
                             in_data[338],
                             in_data[950],
                             in_data[627],
                             in_data[889],
                             in_data[1060],
                             in_data[555]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [63:0] lut_292_table = 64'b1111111011000100111100001100000011110100110001001111011011110100;
    wire [5:0] lut_292_select = {
                             in_data[1068],
                             in_data[987],
                             in_data[2010],
                             in_data[1948],
                             in_data[162],
                             in_data[1043]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [63:0] lut_293_table = 64'b0010001100000001101000110010001100100011000000011011001100110011;
    wire [5:0] lut_293_select = {
                             in_data[1007],
                             in_data[2297],
                             in_data[967],
                             in_data[1940],
                             in_data[906],
                             in_data[1296]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [63:0] lut_294_table = 64'b0000000000000000111011111010111000000000000000001111111110001111;
    wire [5:0] lut_294_select = {
                             in_data[1830],
                             in_data[164],
                             in_data[1945],
                             in_data[2173],
                             in_data[2116],
                             in_data[1288]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [63:0] lut_295_table = 64'b1111000011110000000011000000111001010000000000000000000000000000;
    wire [5:0] lut_295_select = {
                             in_data[361],
                             in_data[1684],
                             in_data[1614],
                             in_data[596],
                             in_data[2138],
                             in_data[1394]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [63:0] lut_296_table = 64'b0000111000001011100011100000100000001111000001010000111000000000;
    wire [5:0] lut_296_select = {
                             in_data[845],
                             in_data[2150],
                             in_data[499],
                             in_data[1871],
                             in_data[129],
                             in_data[81]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [63:0] lut_297_table = 64'b1111111110101010101110110010001011111010101100000000000000000000;
    wire [5:0] lut_297_select = {
                             in_data[1548],
                             in_data[149],
                             in_data[1080],
                             in_data[212],
                             in_data[1084],
                             in_data[185]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [63:0] lut_298_table = 64'b0101000011000000000000000000000011110000110100001110000011000000;
    wire [5:0] lut_298_select = {
                             in_data[1256],
                             in_data[715],
                             in_data[1046],
                             in_data[350],
                             in_data[1542],
                             in_data[1094]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [63:0] lut_299_table = 64'b1111010000001000000001000000000011111101110111011111010100011101;
    wire [5:0] lut_299_select = {
                             in_data[921],
                             in_data[868],
                             in_data[456],
                             in_data[615],
                             in_data[1226],
                             in_data[2002]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [63:0] lut_300_table = 64'b1011001100100010001000110010000000110011001000100010001000000000;
    wire [5:0] lut_300_select = {
                             in_data[484],
                             in_data[169],
                             in_data[2219],
                             in_data[1249],
                             in_data[109],
                             in_data[1885]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [63:0] lut_301_table = 64'b0000110110001111000011011101111111011111111111111111111111111111;
    wire [5:0] lut_301_select = {
                             in_data[1432],
                             in_data[1494],
                             in_data[309],
                             in_data[2231],
                             in_data[1488],
                             in_data[1732]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [63:0] lut_302_table = 64'b1100111111101111111011111111111100000000000011110000000000000000;
    wire [5:0] lut_302_select = {
                             in_data[780],
                             in_data[920],
                             in_data[1627],
                             in_data[1031],
                             in_data[1806],
                             in_data[1604]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [63:0] lut_303_table = 64'b1111111111011100000000001100010011111101111111000000000011010000;
    wire [5:0] lut_303_select = {
                             in_data[2100],
                             in_data[1032],
                             in_data[1950],
                             in_data[154],
                             in_data[1246],
                             in_data[833]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [63:0] lut_304_table = 64'b1010101111101111101010111010101000000011101011110010101110101111;
    wire [5:0] lut_304_select = {
                             in_data[952],
                             in_data[717],
                             in_data[84],
                             in_data[1400],
                             in_data[1327],
                             in_data[1558]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [63:0] lut_305_table = 64'b0000000000100000000000000010001000000000001000100010001000110010;
    wire [5:0] lut_305_select = {
                             in_data[1438],
                             in_data[1821],
                             in_data[1814],
                             in_data[1101],
                             in_data[332],
                             in_data[1967]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [63:0] lut_306_table = 64'b0000000001000100000000000000000001011111111111111101111111111111;
    wire [5:0] lut_306_select = {
                             in_data[1842],
                             in_data[1528],
                             in_data[1216],
                             in_data[1358],
                             in_data[893],
                             in_data[1978]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [63:0] lut_307_table = 64'b0000100000100010010011001111001101001100000100010101110011011111;
    wire [5:0] lut_307_select = {
                             in_data[98],
                             in_data[1497],
                             in_data[2172],
                             in_data[2225],
                             in_data[1556],
                             in_data[2104]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [63:0] lut_308_table = 64'b0100111011111110011100101111111001111110111111101111111111111111;
    wire [5:0] lut_308_select = {
                             in_data[538],
                             in_data[1392],
                             in_data[999],
                             in_data[1415],
                             in_data[919],
                             in_data[2186]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [63:0] lut_309_table = 64'b0111111101011111111110111111111101011111010011111011101011111010;
    wire [5:0] lut_309_select = {
                             in_data[366],
                             in_data[475],
                             in_data[702],
                             in_data[2075],
                             in_data[1239],
                             in_data[68]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [63:0] lut_310_table = 64'b1010111100101010101011101010101011111111101110111111111110111011;
    wire [5:0] lut_310_select = {
                             in_data[1431],
                             in_data[239],
                             in_data[1140],
                             in_data[2020],
                             in_data[132],
                             in_data[853]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [63:0] lut_311_table = 64'b1111111110101111000000100000001000111111111111110000000000000010;
    wire [5:0] lut_311_select = {
                             in_data[1918],
                             in_data[793],
                             in_data[604],
                             in_data[1381],
                             in_data[901],
                             in_data[809]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [63:0] lut_312_table = 64'b0000101010101010000010101010101000000000000000000000000000000000;
    wire [5:0] lut_312_select = {
                             in_data[721],
                             in_data[1322],
                             in_data[1935],
                             in_data[384],
                             in_data[1453],
                             in_data[1673]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [63:0] lut_313_table = 64'b1100000011111111010100010111011101000000111111110000000001010011;
    wire [5:0] lut_313_select = {
                             in_data[1149],
                             in_data[2249],
                             in_data[1880],
                             in_data[2176],
                             in_data[927],
                             in_data[963]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [63:0] lut_314_table = 64'b1000000011111000000000000000000010100000111110000000000010100000;
    wire [5:0] lut_314_select = {
                             in_data[1823],
                             in_data[2194],
                             in_data[1258],
                             in_data[344],
                             in_data[1771],
                             in_data[1766]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [63:0] lut_315_table = 64'b1001111000001000111111111100110000000000000000000000110000001100;
    wire [5:0] lut_315_select = {
                             in_data[167],
                             in_data[1069],
                             in_data[2107],
                             in_data[579],
                             in_data[2137],
                             in_data[677]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [63:0] lut_316_table = 64'b0011011111111111111111111111111100110000111101110010000011110111;
    wire [5:0] lut_316_select = {
                             in_data[537],
                             in_data[737],
                             in_data[834],
                             in_data[1123],
                             in_data[1774],
                             in_data[1440]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [63:0] lut_317_table = 64'b0100110100001100000000000000101001011101010111011100000011111110;
    wire [5:0] lut_317_select = {
                             in_data[1293],
                             in_data[1295],
                             in_data[482],
                             in_data[2261],
                             in_data[954],
                             in_data[543]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [63:0] lut_318_table = 64'b1010100010101110110010001000100010101000101010101000100010001000;
    wire [5:0] lut_318_select = {
                             in_data[1193],
                             in_data[2170],
                             in_data[163],
                             in_data[941],
                             in_data[830],
                             in_data[221]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [63:0] lut_319_table = 64'b1110111010101010110011111111111110101010101010100010101000101011;
    wire [5:0] lut_319_select = {
                             in_data[1275],
                             in_data[589],
                             in_data[298],
                             in_data[2074],
                             in_data[1408],
                             in_data[2096]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [63:0] lut_320_table = 64'b1000000010100000000000001010000011111100101100111111100000110011;
    wire [5:0] lut_320_select = {
                             in_data[377],
                             in_data[923],
                             in_data[1646],
                             in_data[1352],
                             in_data[1388],
                             in_data[4]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [63:0] lut_321_table = 64'b1111111111111111000000000000000011111111111111110000000000000000;
    wire [5:0] lut_321_select = {
                             in_data[296],
                             in_data[479],
                             in_data[2122],
                             in_data[161],
                             in_data[2284],
                             in_data[1265]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [63:0] lut_322_table = 64'b0001000110111001101111111111111100000000000100000011000100110001;
    wire [5:0] lut_322_select = {
                             in_data[2244],
                             in_data[2192],
                             in_data[1026],
                             in_data[1222],
                             in_data[1479],
                             in_data[1891]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [63:0] lut_323_table = 64'b0000000100000001000101110001011100010101000100010101011101010101;
    wire [5:0] lut_323_select = {
                             in_data[1278],
                             in_data[942],
                             in_data[548],
                             in_data[1301],
                             in_data[1397],
                             in_data[1146]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [63:0] lut_324_table = 64'b0101010101010111111111101101111001010101010101110101000001010000;
    wire [5:0] lut_324_select = {
                             in_data[8],
                             in_data[307],
                             in_data[2287],
                             in_data[412],
                             in_data[1653],
                             in_data[1206]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [63:0] lut_325_table = 64'b0110011001100010011001110110011111111110111001000110111101000110;
    wire [5:0] lut_325_select = {
                             in_data[666],
                             in_data[815],
                             in_data[1477],
                             in_data[2001],
                             in_data[1349],
                             in_data[770]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [63:0] lut_326_table = 64'b0000100010111010000110011111101111010000111100011111000111110001;
    wire [5:0] lut_326_select = {
                             in_data[1701],
                             in_data[1390],
                             in_data[76],
                             in_data[1472],
                             in_data[1547],
                             in_data[1841]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [63:0] lut_327_table = 64'b1111010110110000111111011111000011111101101100011111110110111001;
    wire [5:0] lut_327_select = {
                             in_data[1616],
                             in_data[408],
                             in_data[1041],
                             in_data[623],
                             in_data[752],
                             in_data[2187]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [63:0] lut_328_table = 64'b0010000100110011000000000111011100100000101100110000000000110011;
    wire [5:0] lut_328_select = {
                             in_data[2112],
                             in_data[536],
                             in_data[1803],
                             in_data[2127],
                             in_data[513],
                             in_data[147]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [63:0] lut_329_table = 64'b0000001100010111001101110101011100001000010001010000110101010101;
    wire [5:0] lut_329_select = {
                             in_data[2049],
                             in_data[763],
                             in_data[1332],
                             in_data[358],
                             in_data[678],
                             in_data[1852]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [63:0] lut_330_table = 64'b0101111111010101110101011101010111110000110100001111000011010000;
    wire [5:0] lut_330_select = {
                             in_data[570],
                             in_data[1822],
                             in_data[2184],
                             in_data[565],
                             in_data[551],
                             in_data[1436]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [63:0] lut_331_table = 64'b1100110010000000110011001000000010001000000000001000100000000000;
    wire [5:0] lut_331_select = {
                             in_data[2153],
                             in_data[1331],
                             in_data[1052],
                             in_data[769],
                             in_data[468],
                             in_data[2136]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [63:0] lut_332_table = 64'b0011011100000000011111110010000000000111000000010000111100000001;
    wire [5:0] lut_332_select = {
                             in_data[341],
                             in_data[1124],
                             in_data[2274],
                             in_data[530],
                             in_data[1845],
                             in_data[587]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [63:0] lut_333_table = 64'b0101010100001101110111010101110101010101000101010111010101010101;
    wire [5:0] lut_333_select = {
                             in_data[52],
                             in_data[598],
                             in_data[1437],
                             in_data[1045],
                             in_data[112],
                             in_data[1200]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [63:0] lut_334_table = 64'b0001000100010111000100010001011100010001111111110001000011111111;
    wire [5:0] lut_334_select = {
                             in_data[312],
                             in_data[480],
                             in_data[713],
                             in_data[1742],
                             in_data[1815],
                             in_data[49]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [63:0] lut_335_table = 64'b0101000011110111011100110111001101110001111100110111001101110011;
    wire [5:0] lut_335_select = {
                             in_data[1180],
                             in_data[676],
                             in_data[2212],
                             in_data[1867],
                             in_data[1717],
                             in_data[447]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [63:0] lut_336_table = 64'b0010000000100000001000000000000011110000111100001011000000010000;
    wire [5:0] lut_336_select = {
                             in_data[1763],
                             in_data[1539],
                             in_data[1441],
                             in_data[636],
                             in_data[1082],
                             in_data[723]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [63:0] lut_337_table = 64'b0000101000001010000111110000101100001010001010100001000101010111;
    wire [5:0] lut_337_select = {
                             in_data[683],
                             in_data[1809],
                             in_data[1743],
                             in_data[1892],
                             in_data[2018],
                             in_data[1459]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [63:0] lut_338_table = 64'b1111111111111111101100101011001111111111111111111011000010110011;
    wire [5:0] lut_338_select = {
                             in_data[201],
                             in_data[2234],
                             in_data[918],
                             in_data[385],
                             in_data[1345],
                             in_data[1734]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [63:0] lut_339_table = 64'b0000001101001111010011110101011100000010000000110101101101010011;
    wire [5:0] lut_339_select = {
                             in_data[2110],
                             in_data[2163],
                             in_data[1366],
                             in_data[992],
                             in_data[907],
                             in_data[1071]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [63:0] lut_340_table = 64'b1110111011111110110011001100111011101010111111101100000011000000;
    wire [5:0] lut_340_select = {
                             in_data[508],
                             in_data[1030],
                             in_data[268],
                             in_data[2197],
                             in_data[991],
                             in_data[2247]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [63:0] lut_341_table = 64'b1000111000001010101011111111011110000000000000000100000011110000;
    wire [5:0] lut_341_select = {
                             in_data[1173],
                             in_data[265],
                             in_data[1862],
                             in_data[1009],
                             in_data[2199],
                             in_data[944]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [63:0] lut_342_table = 64'b1101010101000001110000000000000111111111010101111100010101000101;
    wire [5:0] lut_342_select = {
                             in_data[253],
                             in_data[2237],
                             in_data[2168],
                             in_data[392],
                             in_data[1356],
                             in_data[1230]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [63:0] lut_343_table = 64'b1110000011101010001000001100010010110010111111110000000010100000;
    wire [5:0] lut_343_select = {
                             in_data[808],
                             in_data[583],
                             in_data[1678],
                             in_data[695],
                             in_data[191],
                             in_data[811]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [63:0] lut_344_table = 64'b0000010000001100000111110001111110101100101111001111111100011101;
    wire [5:0] lut_344_select = {
                             in_data[1103],
                             in_data[1733],
                             in_data[54],
                             in_data[751],
                             in_data[151],
                             in_data[2256]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [63:0] lut_345_table = 64'b1111001111111011001100000000000000100000001000000000000000000000;
    wire [5:0] lut_345_select = {
                             in_data[1668],
                             in_data[339],
                             in_data[1554],
                             in_data[1442],
                             in_data[1937],
                             in_data[1445]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [63:0] lut_346_table = 64'b1110111100001110111111110000111101000110000000000100111100000101;
    wire [5:0] lut_346_select = {
                             in_data[155],
                             in_data[710],
                             in_data[355],
                             in_data[254],
                             in_data[224],
                             in_data[1747]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [63:0] lut_347_table = 64'b1111001100110000111100110011001000110001001100001111001100110010;
    wire [5:0] lut_347_select = {
                             in_data[134],
                             in_data[381],
                             in_data[1023],
                             in_data[122],
                             in_data[1591],
                             in_data[1648]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [63:0] lut_348_table = 64'b1111111011111110110011001111111011101100110011001100000011001100;
    wire [5:0] lut_348_select = {
                             in_data[1471],
                             in_data[1714],
                             in_data[787],
                             in_data[909],
                             in_data[524],
                             in_data[249]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [63:0] lut_349_table = 64'b1111010011101101011100000000010011111110101011001111000000000000;
    wire [5:0] lut_349_select = {
                             in_data[759],
                             in_data[1920],
                             in_data[1402],
                             in_data[1998],
                             in_data[1761],
                             in_data[1053]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [63:0] lut_350_table = 64'b0101010011111111111111111111111100000000000000010101110100000011;
    wire [5:0] lut_350_select = {
                             in_data[2190],
                             in_data[1398],
                             in_data[1569],
                             in_data[2240],
                             in_data[1153],
                             in_data[2062]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [63:0] lut_351_table = 64'b0000000001010000010000001101010000000000010101010000000011010101;
    wire [5:0] lut_351_select = {
                             in_data[995],
                             in_data[1414],
                             in_data[2250],
                             in_data[1245],
                             in_data[739],
                             in_data[884]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [63:0] lut_352_table = 64'b1111110011111111110010001111000011101000111111111100100011101010;
    wire [5:0] lut_352_select = {
                             in_data[1166],
                             in_data[60],
                             in_data[783],
                             in_data[1762],
                             in_data[772],
                             in_data[882]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [63:0] lut_353_table = 64'b0010101000101110000010001111111110101010101010100011101011111111;
    wire [5:0] lut_353_select = {
                             in_data[754],
                             in_data[46],
                             in_data[386],
                             in_data[1644],
                             in_data[1422],
                             in_data[1439]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [63:0] lut_354_table = 64'b0101010100000000010101010001000100010001000000000001000100000000;
    wire [5:0] lut_354_select = {
                             in_data[1658],
                             in_data[554],
                             in_data[973],
                             in_data[730],
                             in_data[1399],
                             in_data[514]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [63:0] lut_355_table = 64'b1110110011111100101011001110110011111100111111001111100011111100;
    wire [5:0] lut_355_select = {
                             in_data[1603],
                             in_data[1446],
                             in_data[1059],
                             in_data[248],
                             in_data[888],
                             in_data[571]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [63:0] lut_356_table = 64'b0000100000000010101011101010111011101111111011110010111111101111;
    wire [5:0] lut_356_select = {
                             in_data[1487],
                             in_data[291],
                             in_data[1520],
                             in_data[1129],
                             in_data[1120],
                             in_data[669]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [63:0] lut_357_table = 64'b0101110100000000110111110000000000000000000000000100010001010101;
    wire [5:0] lut_357_select = {
                             in_data[1605],
                             in_data[1412],
                             in_data[660],
                             in_data[1557],
                             in_data[40],
                             in_data[1308]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [63:0] lut_358_table = 64'b1110111111101111101011111000110100000000000001001000110010000100;
    wire [5:0] lut_358_select = {
                             in_data[2071],
                             in_data[512],
                             in_data[504],
                             in_data[1719],
                             in_data[1915],
                             in_data[1608]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [63:0] lut_359_table = 64'b0101010101010001010100000101000011110101111101010111010101110101;
    wire [5:0] lut_359_select = {
                             in_data[1578],
                             in_data[94],
                             in_data[1168],
                             in_data[1595],
                             in_data[854],
                             in_data[399]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [63:0] lut_360_table = 64'b0101010101000000010001000000000011111111111111111101010111111100;
    wire [5:0] lut_360_select = {
                             in_data[2011],
                             in_data[443],
                             in_data[517],
                             in_data[2270],
                             in_data[1857],
                             in_data[1022]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [63:0] lut_361_table = 64'b0011011100110001011111110001000101110111011101010111111100110101;
    wire [5:0] lut_361_select = {
                             in_data[646],
                             in_data[2233],
                             in_data[857],
                             in_data[1698],
                             in_data[819],
                             in_data[1795]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [63:0] lut_362_table = 64'b0100010000000000110011011100110101000101010001001100110111001101;
    wire [5:0] lut_362_select = {
                             in_data[1516],
                             in_data[994],
                             in_data[329],
                             in_data[2088],
                             in_data[1875],
                             in_data[1586]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [63:0] lut_363_table = 64'b1111111101110011001110110000000011111111111111110011011100010001;
    wire [5:0] lut_363_select = {
                             in_data[292],
                             in_data[204],
                             in_data[334],
                             in_data[523],
                             in_data[980],
                             in_data[1599]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [63:0] lut_364_table = 64'b1111111101001101000111110000010111001111000010001111111100000000;
    wire [5:0] lut_364_select = {
                             in_data[29],
                             in_data[561],
                             in_data[1463],
                             in_data[1170],
                             in_data[2139],
                             in_data[617]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [63:0] lut_365_table = 64'b1111000011000000011100100011000001110010010100000111001101110011;
    wire [5:0] lut_365_select = {
                             in_data[67],
                             in_data[1252],
                             in_data[984],
                             in_data[1027],
                             in_data[336],
                             in_data[186]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [63:0] lut_366_table = 64'b0000101000100011001000100010001110111111111111111111001111111111;
    wire [5:0] lut_366_select = {
                             in_data[1654],
                             in_data[1941],
                             in_data[1567],
                             in_data[1391],
                             in_data[409],
                             in_data[250]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [63:0] lut_367_table = 64'b1101111111011100110111111101110011011111111111110100111111011100;
    wire [5:0] lut_367_select = {
                             in_data[1135],
                             in_data[2014],
                             in_data[765],
                             in_data[2045],
                             in_data[2008],
                             in_data[1923]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [63:0] lut_368_table = 64'b1100110001001100010011000000110011001100110010001100110010001000;
    wire [5:0] lut_368_select = {
                             in_data[2039],
                             in_data[859],
                             in_data[1297],
                             in_data[13],
                             in_data[1346],
                             in_data[2147]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [63:0] lut_369_table = 64'b0111001101010001111110110101001111110111011100011100000001010001;
    wire [5:0] lut_369_select = {
                             in_data[625],
                             in_data[2232],
                             in_data[1443],
                             in_data[2103],
                             in_data[1002],
                             in_data[2245]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [63:0] lut_370_table = 64'b1111111111111111000000110000000011111111111111111011101111111011;
    wire [5:0] lut_370_select = {
                             in_data[2175],
                             in_data[1794],
                             in_data[2142],
                             in_data[2081],
                             in_data[333],
                             in_data[1204]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [63:0] lut_371_table = 64'b0100000001000000110101001100010001000000000000001111110011000100;
    wire [5:0] lut_371_select = {
                             in_data[281],
                             in_data[1385],
                             in_data[1161],
                             in_data[469],
                             in_data[2217],
                             in_data[969]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [63:0] lut_372_table = 64'b0001000000011011011100010001111100000000000000000101000000000001;
    wire [5:0] lut_372_select = {
                             in_data[319],
                             in_data[1526],
                             in_data[1197],
                             in_data[934],
                             in_data[246],
                             in_data[983]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [63:0] lut_373_table = 64'b0111000001110101001100110111011101110011111101110011001111111111;
    wire [5:0] lut_373_select = {
                             in_data[200],
                             in_data[692],
                             in_data[2288],
                             in_data[465],
                             in_data[121],
                             in_data[564]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [63:0] lut_374_table = 64'b1111000001010000000001000000110011111110111111101100111010001100;
    wire [5:0] lut_374_select = {
                             in_data[502],
                             in_data[729],
                             in_data[1713],
                             in_data[1607],
                             in_data[1454],
                             in_data[2134]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [63:0] lut_375_table = 64'b0111101000001011000000000000101011111111110111110100100010001100;
    wire [5:0] lut_375_select = {
                             in_data[337],
                             in_data[431],
                             in_data[400],
                             in_data[903],
                             in_data[243],
                             in_data[1514]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [63:0] lut_376_table = 64'b1111011111111111111100001111000010101010100010101010101000000010;
    wire [5:0] lut_376_select = {
                             in_data[1921],
                             in_data[1635],
                             in_data[2182],
                             in_data[1898],
                             in_data[1070],
                             in_data[419]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [63:0] lut_377_table = 64'b1111111000111010101111000000100011111100000111111101110000001100;
    wire [5:0] lut_377_select = {
                             in_data[1138],
                             in_data[978],
                             in_data[1421],
                             in_data[90],
                             in_data[535],
                             in_data[779]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [63:0] lut_378_table = 64'b1010101010101010101010001000100011101110111011101010111010001000;
    wire [5:0] lut_378_select = {
                             in_data[2277],
                             in_data[861],
                             in_data[158],
                             in_data[467],
                             in_data[1980],
                             in_data[2258]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [63:0] lut_379_table = 64'b0010001000000000111111110010101000100010000000000011001000100000;
    wire [5:0] lut_379_select = {
                             in_data[133],
                             in_data[1100],
                             in_data[829],
                             in_data[1835],
                             in_data[476],
                             in_data[2296]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [63:0] lut_380_table = 64'b0000010000001100010011001101110000000000000000000100110001011100;
    wire [5:0] lut_380_select = {
                             in_data[2098],
                             in_data[225],
                             in_data[711],
                             in_data[335],
                             in_data[1355],
                             in_data[814]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [63:0] lut_381_table = 64'b1111111100001101111111110100110111111111110111111111111111011101;
    wire [5:0] lut_381_select = {
                             in_data[1110],
                             in_data[803],
                             in_data[1901],
                             in_data[451],
                             in_data[1096],
                             in_data[1189]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [63:0] lut_382_table = 64'b1010111110001111101010101000101010000100100011011010000010000000;
    wire [5:0] lut_382_select = {
                             in_data[503],
                             in_data[2114],
                             in_data[1666],
                             in_data[188],
                             in_data[790],
                             in_data[1824]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [63:0] lut_383_table = 64'b1100010000000000110111001111110111010100111111011101110011111101;
    wire [5:0] lut_383_select = {
                             in_data[198],
                             in_data[1729],
                             in_data[1426],
                             in_data[1805],
                             in_data[2145],
                             in_data[1688]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub2
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        383:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [         63:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub2_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub2_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub2_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [383:0]  in_data,
            output wire [63:0]  out_data
        );
    
    
    // LUT : 0
    wire [63:0] lut_0_table = 64'b0001111100000101111111111101111100000000000000000001011100010111;
    wire [5:0] lut_0_select = {
                             in_data[111],
                             in_data[82],
                             in_data[280],
                             in_data[316],
                             in_data[302],
                             in_data[8]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [63:0] lut_1_table = 64'b1000100000001100000000000000101011111111000011101010101000001110;
    wire [5:0] lut_1_select = {
                             in_data[20],
                             in_data[289],
                             in_data[203],
                             in_data[344],
                             in_data[191],
                             in_data[73]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [63:0] lut_2_table = 64'b1110000011101100111111101110111110000000101000001110100010101010;
    wire [5:0] lut_2_select = {
                             in_data[310],
                             in_data[148],
                             in_data[47],
                             in_data[10],
                             in_data[278],
                             in_data[71]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [63:0] lut_3_table = 64'b0000000000000001000001010101011100000111011111110001111111111111;
    wire [5:0] lut_3_select = {
                             in_data[330],
                             in_data[120],
                             in_data[98],
                             in_data[178],
                             in_data[44],
                             in_data[133]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [63:0] lut_4_table = 64'b1111110111011100110101010100000011000100110001001100010000000000;
    wire [5:0] lut_4_select = {
                             in_data[132],
                             in_data[234],
                             in_data[48],
                             in_data[129],
                             in_data[259],
                             in_data[334]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [63:0] lut_5_table = 64'b1000111010001000111011101111111100001000000010001000111011101110;
    wire [5:0] lut_5_select = {
                             in_data[0],
                             in_data[65],
                             in_data[30],
                             in_data[193],
                             in_data[298],
                             in_data[41]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [63:0] lut_6_table = 64'b1101010011010100010000000100000011111101110111001101010111000100;
    wire [5:0] lut_6_select = {
                             in_data[206],
                             in_data[359],
                             in_data[347],
                             in_data[40],
                             in_data[135],
                             in_data[205]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [63:0] lut_7_table = 64'b0000110000001100100011101100111111001000110011001100110011001111;
    wire [5:0] lut_7_select = {
                             in_data[338],
                             in_data[341],
                             in_data[61],
                             in_data[254],
                             in_data[320],
                             in_data[275]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [63:0] lut_8_table = 64'b1111111111011101110101000000000011111100110000001101010000000000;
    wire [5:0] lut_8_select = {
                             in_data[200],
                             in_data[101],
                             in_data[371],
                             in_data[274],
                             in_data[78],
                             in_data[329]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [63:0] lut_9_table = 64'b0000001000000000100000100010011110101011101011111010001000101111;
    wire [5:0] lut_9_select = {
                             in_data[378],
                             in_data[322],
                             in_data[265],
                             in_data[327],
                             in_data[141],
                             in_data[355]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [63:0] lut_10_table = 64'b1111111111001101110011000000000011111111110111111101110111001101;
    wire [5:0] lut_10_select = {
                             in_data[218],
                             in_data[235],
                             in_data[252],
                             in_data[37],
                             in_data[36],
                             in_data[296]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [63:0] lut_11_table = 64'b0100010101001100010011000100110101011101110111011100110111111111;
    wire [5:0] lut_11_select = {
                             in_data[125],
                             in_data[159],
                             in_data[124],
                             in_data[32],
                             in_data[53],
                             in_data[224]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [63:0] lut_12_table = 64'b0000110000000000110111000000110001011111000011001101111111011100;
    wire [5:0] lut_12_select = {
                             in_data[123],
                             in_data[147],
                             in_data[340],
                             in_data[115],
                             in_data[171],
                             in_data[369]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [63:0] lut_13_table = 64'b0001000100010000011101010111000001010001000100001111011111110000;
    wire [5:0] lut_13_select = {
                             in_data[181],
                             in_data[376],
                             in_data[263],
                             in_data[168],
                             in_data[128],
                             in_data[232]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [63:0] lut_14_table = 64'b1101110111001100010001010000000011011111110111010101110100001100;
    wire [5:0] lut_14_select = {
                             in_data[293],
                             in_data[276],
                             in_data[352],
                             in_data[104],
                             in_data[19],
                             in_data[94]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [63:0] lut_15_table = 64'b0011000001110111011100010111010100000000000100010001000101110101;
    wire [5:0] lut_15_select = {
                             in_data[144],
                             in_data[79],
                             in_data[267],
                             in_data[272],
                             in_data[317],
                             in_data[112]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [63:0] lut_16_table = 64'b0100010011110101110111001111111100000000010101000100000011110101;
    wire [5:0] lut_16_select = {
                             in_data[353],
                             in_data[116],
                             in_data[337],
                             in_data[58],
                             in_data[97],
                             in_data[368]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [63:0] lut_17_table = 64'b0101000011110111000100001010000001110001111111110111000011111011;
    wire [5:0] lut_17_select = {
                             in_data[304],
                             in_data[221],
                             in_data[182],
                             in_data[34],
                             in_data[319],
                             in_data[77]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [63:0] lut_18_table = 64'b0000111001001000000010101110111010001110000010000000000000000000;
    wire [5:0] lut_18_select = {
                             in_data[152],
                             in_data[216],
                             in_data[33],
                             in_data[167],
                             in_data[374],
                             in_data[339]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [63:0] lut_19_table = 64'b0110111111111111111111111111111100000010001010100010101110111111;
    wire [5:0] lut_19_select = {
                             in_data[74],
                             in_data[45],
                             in_data[315],
                             in_data[4],
                             in_data[365],
                             in_data[166]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [63:0] lut_20_table = 64'b0010001110111111001000101010101110111011101111110010101110101111;
    wire [5:0] lut_20_select = {
                             in_data[64],
                             in_data[266],
                             in_data[262],
                             in_data[312],
                             in_data[172],
                             in_data[21]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [63:0] lut_21_table = 64'b0000000011110101100000001111010110110001111101110001000011110111;
    wire [5:0] lut_21_select = {
                             in_data[54],
                             in_data[311],
                             in_data[211],
                             in_data[51],
                             in_data[26],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [63:0] lut_22_table = 64'b1011000011110010101100101111001100100000001100000010000000110000;
    wire [5:0] lut_22_select = {
                             in_data[43],
                             in_data[107],
                             in_data[1],
                             in_data[52],
                             in_data[332],
                             in_data[118]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [63:0] lut_23_table = 64'b0001000101010111000000000000000111111111111111111000101111111111;
    wire [5:0] lut_23_select = {
                             in_data[202],
                             in_data[188],
                             in_data[195],
                             in_data[335],
                             in_data[49],
                             in_data[35]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [63:0] lut_24_table = 64'b1111111011111101111010100000110011111000100000001110100000000000;
    wire [5:0] lut_24_select = {
                             in_data[17],
                             in_data[155],
                             in_data[270],
                             in_data[241],
                             in_data[149],
                             in_data[269]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [63:0] lut_25_table = 64'b0000010001000100010001001111111101000101010101010101110111111111;
    wire [5:0] lut_25_select = {
                             in_data[63],
                             in_data[69],
                             in_data[248],
                             in_data[142],
                             in_data[176],
                             in_data[357]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [63:0] lut_26_table = 64'b0001011100000001011111110011001100010001000000000001011100000001;
    wire [5:0] lut_26_select = {
                             in_data[361],
                             in_data[236],
                             in_data[324],
                             in_data[11],
                             in_data[179],
                             in_data[131]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [63:0] lut_27_table = 64'b0011111111111111000101110111111100000000000101110000000100010111;
    wire [5:0] lut_27_select = {
                             in_data[16],
                             in_data[164],
                             in_data[256],
                             in_data[223],
                             in_data[122],
                             in_data[86]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [63:0] lut_28_table = 64'b0000001000100010001010111011101100100010101110111011101111111111;
    wire [5:0] lut_28_select = {
                             in_data[80],
                             in_data[346],
                             in_data[84],
                             in_data[244],
                             in_data[2],
                             in_data[283]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [63:0] lut_29_table = 64'b1000100110001000000010010000100011011111110011111000100110001000;
    wire [5:0] lut_29_select = {
                             in_data[264],
                             in_data[130],
                             in_data[186],
                             in_data[249],
                             in_data[42],
                             in_data[331]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [63:0] lut_30_table = 64'b1110110011101111101010001110110010001000111011111010100010101000;
    wire [5:0] lut_30_select = {
                             in_data[286],
                             in_data[99],
                             in_data[284],
                             in_data[333],
                             in_data[151],
                             in_data[321]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [63:0] lut_31_table = 64'b0001000100111111001101110111111100000000001100010001000100110111;
    wire [5:0] lut_31_select = {
                             in_data[228],
                             in_data[67],
                             in_data[160],
                             in_data[3],
                             in_data[189],
                             in_data[243]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [63:0] lut_32_table = 64'b1111101011101111101010101000111111111111111111111010101011111111;
    wire [5:0] lut_32_select = {
                             in_data[60],
                             in_data[62],
                             in_data[294],
                             in_data[198],
                             in_data[229],
                             in_data[309]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [63:0] lut_33_table = 64'b0000000000000010001110110000101000111011000000101111111100111011;
    wire [5:0] lut_33_select = {
                             in_data[214],
                             in_data[100],
                             in_data[318],
                             in_data[207],
                             in_data[204],
                             in_data[39]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [63:0] lut_34_table = 64'b0000000000110010001000001011101100110010101110111011001011111011;
    wire [5:0] lut_34_select = {
                             in_data[292],
                             in_data[279],
                             in_data[76],
                             in_data[81],
                             in_data[197],
                             in_data[113]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [63:0] lut_35_table = 64'b0000010001001111010011000101011100001100010111110100110111011111;
    wire [5:0] lut_35_select = {
                             in_data[190],
                             in_data[14],
                             in_data[209],
                             in_data[177],
                             in_data[92],
                             in_data[314]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [63:0] lut_36_table = 64'b1111001101110001111101110111001101110001000100000111000100010001;
    wire [5:0] lut_36_select = {
                             in_data[240],
                             in_data[27],
                             in_data[370],
                             in_data[367],
                             in_data[287],
                             in_data[273]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [63:0] lut_37_table = 64'b0101010111111111000000001111110101110001111101110101000111110111;
    wire [5:0] lut_37_select = {
                             in_data[22],
                             in_data[46],
                             in_data[381],
                             in_data[323],
                             in_data[362],
                             in_data[134]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [63:0] lut_38_table = 64'b0111001111111111001100011111011100010000011101110000000000010001;
    wire [5:0] lut_38_select = {
                             in_data[119],
                             in_data[251],
                             in_data[169],
                             in_data[183],
                             in_data[162],
                             in_data[108]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [63:0] lut_39_table = 64'b1000111011101110101011101110111100000000100011001000100010101110;
    wire [5:0] lut_39_select = {
                             in_data[253],
                             in_data[215],
                             in_data[114],
                             in_data[28],
                             in_data[336],
                             in_data[328]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [63:0] lut_40_table = 64'b0000111010101111000000100000101110001110111111110010101110101111;
    wire [5:0] lut_40_select = {
                             in_data[364],
                             in_data[173],
                             in_data[326],
                             in_data[127],
                             in_data[5],
                             in_data[25]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [63:0] lut_41_table = 64'b1100111100001101010011010000000011011111110011111101111100001101;
    wire [5:0] lut_41_select = {
                             in_data[210],
                             in_data[68],
                             in_data[225],
                             in_data[12],
                             in_data[345],
                             in_data[174]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [63:0] lut_42_table = 64'b1011001111111011101000001111100100110000111100100010000010110000;
    wire [5:0] lut_42_select = {
                             in_data[238],
                             in_data[139],
                             in_data[93],
                             in_data[380],
                             in_data[89],
                             in_data[379]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [63:0] lut_43_table = 64'b0000010101010001000000010011001101011111111111110001011100111111;
    wire [5:0] lut_43_select = {
                             in_data[271],
                             in_data[138],
                             in_data[105],
                             in_data[307],
                             in_data[66],
                             in_data[91]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [63:0] lut_44_table = 64'b0101100001001000000000000000000011111101110111011000110010011000;
    wire [5:0] lut_44_select = {
                             in_data[150],
                             in_data[90],
                             in_data[301],
                             in_data[233],
                             in_data[95],
                             in_data[137]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [63:0] lut_45_table = 64'b1010111110001110000010000000100011111111101011111100111110001110;
    wire [5:0] lut_45_select = {
                             in_data[373],
                             in_data[59],
                             in_data[145],
                             in_data[308],
                             in_data[299],
                             in_data[13]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [63:0] lut_46_table = 64'b1000100011101110111010101111111110001100110011101110110011101111;
    wire [5:0] lut_46_select = {
                             in_data[383],
                             in_data[170],
                             in_data[250],
                             in_data[354],
                             in_data[261],
                             in_data[121]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [63:0] lut_47_table = 64'b1111111111111010111110101011000011111010111110001011000010000000;
    wire [5:0] lut_47_select = {
                             in_data[297],
                             in_data[70],
                             in_data[285],
                             in_data[288],
                             in_data[180],
                             in_data[83]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [63:0] lut_48_table = 64'b1100111111001101111011111100111100001110010011011100111011001111;
    wire [5:0] lut_48_select = {
                             in_data[55],
                             in_data[184],
                             in_data[117],
                             in_data[303],
                             in_data[245],
                             in_data[349]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [63:0] lut_49_table = 64'b1111111011111111111110001101111011011101110111110100000001001100;
    wire [5:0] lut_49_select = {
                             in_data[246],
                             in_data[375],
                             in_data[163],
                             in_data[50],
                             in_data[140],
                             in_data[56]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [63:0] lut_50_table = 64'b1111001101010000111100110111000001110101000100011111111111110001;
    wire [5:0] lut_50_select = {
                             in_data[306],
                             in_data[363],
                             in_data[277],
                             in_data[268],
                             in_data[358],
                             in_data[109]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [63:0] lut_51_table = 64'b1011101010100000101000000010000011111111111110111111111110100000;
    wire [5:0] lut_51_select = {
                             in_data[219],
                             in_data[213],
                             in_data[305],
                             in_data[9],
                             in_data[143],
                             in_data[199]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [63:0] lut_52_table = 64'b0010001010101111001000100010101100100010001111110010001000101011;
    wire [5:0] lut_52_select = {
                             in_data[165],
                             in_data[154],
                             in_data[126],
                             in_data[87],
                             in_data[31],
                             in_data[342]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [63:0] lut_53_table = 64'b1110100010100000111100001111000011111010111010001111111011111010;
    wire [5:0] lut_53_select = {
                             in_data[7],
                             in_data[153],
                             in_data[300],
                             in_data[212],
                             in_data[281],
                             in_data[192]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [63:0] lut_54_table = 64'b0111011100010101000101110000000111111111010111110111111100010111;
    wire [5:0] lut_54_select = {
                             in_data[23],
                             in_data[313],
                             in_data[239],
                             in_data[6],
                             in_data[110],
                             in_data[29]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [63:0] lut_55_table = 64'b0000101000001010001010111010101100001010100011100010101110101111;
    wire [5:0] lut_55_select = {
                             in_data[255],
                             in_data[15],
                             in_data[227],
                             in_data[85],
                             in_data[18],
                             in_data[196]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [63:0] lut_56_table = 64'b1111000011111101000000001101000011111101111111111111000011111101;
    wire [5:0] lut_56_select = {
                             in_data[38],
                             in_data[217],
                             in_data[106],
                             in_data[103],
                             in_data[57],
                             in_data[24]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [63:0] lut_57_table = 64'b0100111111111111010101011101110111011111111111110101110111011111;
    wire [5:0] lut_57_select = {
                             in_data[366],
                             in_data[146],
                             in_data[156],
                             in_data[242],
                             in_data[377],
                             in_data[257]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [63:0] lut_58_table = 64'b1111011101110001000100000000000011111111111101010111000000010000;
    wire [5:0] lut_58_select = {
                             in_data[185],
                             in_data[158],
                             in_data[350],
                             in_data[343],
                             in_data[325],
                             in_data[88]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [63:0] lut_59_table = 64'b0010101000101111101111111111111100000000000010000010101011111111;
    wire [5:0] lut_59_select = {
                             in_data[72],
                             in_data[295],
                             in_data[258],
                             in_data[187],
                             in_data[348],
                             in_data[372]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [63:0] lut_60_table = 64'b1100000011111100000000001100000011011100111111001100000011101100;
    wire [5:0] lut_60_select = {
                             in_data[220],
                             in_data[75],
                             in_data[356],
                             in_data[351],
                             in_data[231],
                             in_data[291]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [63:0] lut_61_table = 64'b1000101010001110100010100000100011111111110011101110111101001100;
    wire [5:0] lut_61_select = {
                             in_data[194],
                             in_data[290],
                             in_data[96],
                             in_data[247],
                             in_data[136],
                             in_data[237]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [63:0] lut_62_table = 64'b0111001011111111011100110111111100000010011101110000000000010011;
    wire [5:0] lut_62_select = {
                             in_data[282],
                             in_data[222],
                             in_data[161],
                             in_data[360],
                             in_data[260],
                             in_data[201]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [63:0] lut_63_table = 64'b1111111111101111111011111000110011101111100011101000111000000000;
    wire [5:0] lut_63_select = {
                             in_data[226],
                             in_data[230],
                             in_data[102],
                             in_data[175],
                             in_data[382],
                             in_data[157]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub3
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [         63:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        359:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub3_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub3_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub3_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [63:0]  in_data,
            output wire [359:0]  out_data
        );
    
    
    // LUT : 0
    wire [63:0] lut_0_table = 64'b0011101000111011101100001011101000111101111111110011000011110100;
    wire [5:0] lut_0_select = {
                             in_data[33],
                             in_data[52],
                             in_data[32],
                             in_data[27],
                             in_data[17],
                             in_data[8]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [63:0] lut_1_table = 64'b1111111111110000111111110101000011111111001000001111111100000000;
    wire [5:0] lut_1_select = {
                             in_data[20],
                             in_data[53],
                             in_data[14],
                             in_data[26],
                             in_data[25],
                             in_data[51]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [63:0] lut_2_table = 64'b1111101110111010101010101011101000110000101110100011001010111010;
    wire [5:0] lut_2_select = {
                             in_data[57],
                             in_data[63],
                             in_data[47],
                             in_data[10],
                             in_data[3],
                             in_data[24]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [63:0] lut_3_table = 64'b0000101010011010000010101000101000001010111110100000101000001000;
    wire [5:0] lut_3_select = {
                             in_data[62],
                             in_data[21],
                             in_data[58],
                             in_data[22],
                             in_data[44],
                             in_data[19]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [63:0] lut_4_table = 64'b1111001001010000111101111101010101000000010100001101010011010101;
    wire [5:0] lut_4_select = {
                             in_data[45],
                             in_data[31],
                             in_data[48],
                             in_data[9],
                             in_data[7],
                             in_data[15]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [63:0] lut_5_table = 64'b0101010101000100110101011100010001010101010001000101010101010100;
    wire [5:0] lut_5_select = {
                             in_data[0],
                             in_data[28],
                             in_data[30],
                             in_data[34],
                             in_data[2],
                             in_data[41]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [63:0] lut_6_table = 64'b1111111100111011000111110000000010111111001000100011111100000000;
    wire [5:0] lut_6_select = {
                             in_data[18],
                             in_data[54],
                             in_data[35],
                             in_data[40],
                             in_data[1],
                             in_data[60]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [63:0] lut_7_table = 64'b0010000000000000111011110000110100100010000000001110111000001101;
    wire [5:0] lut_7_select = {
                             in_data[46],
                             in_data[38],
                             in_data[61],
                             in_data[42],
                             in_data[6],
                             in_data[4]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [63:0] lut_8_table = 64'b1110101010000000111011101110101010101000000000001110101010000000;
    wire [5:0] lut_8_select = {
                             in_data[13],
                             in_data[29],
                             in_data[39],
                             in_data[59],
                             in_data[11],
                             in_data[23]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [63:0] lut_9_table = 64'b1010101010101010111011101010100010001100100010001111111111111100;
    wire [5:0] lut_9_select = {
                             in_data[43],
                             in_data[12],
                             in_data[49],
                             in_data[55],
                             in_data[56],
                             in_data[5]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [63:0] lut_10_table = 64'b0101010111000100010100000101000011110111011111110111010101110101;
    wire [5:0] lut_10_select = {
                             in_data[58],
                             in_data[9],
                             in_data[16],
                             in_data[37],
                             in_data[36],
                             in_data[50]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [63:0] lut_11_table = 64'b1010101110101010101000101000000010111011101110111111101111110010;
    wire [5:0] lut_11_select = {
                             in_data[28],
                             in_data[27],
                             in_data[51],
                             in_data[26],
                             in_data[11],
                             in_data[6]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [63:0] lut_12_table = 64'b0011111111111111000000011111111100000011000100010000000010010011;
    wire [5:0] lut_12_select = {
                             in_data[5],
                             in_data[45],
                             in_data[25],
                             in_data[55],
                             in_data[10],
                             in_data[61]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [63:0] lut_13_table = 64'b0010000010100000101100101111101000100000101011101011001011111111;
    wire [5:0] lut_13_select = {
                             in_data[2],
                             in_data[22],
                             in_data[59],
                             in_data[43],
                             in_data[60],
                             in_data[24]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [63:0] lut_14_table = 64'b1111111101011111011111110001111101010101000011000001010100000000;
    wire [5:0] lut_14_select = {
                             in_data[21],
                             in_data[35],
                             in_data[3],
                             in_data[32],
                             in_data[1],
                             in_data[20]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [63:0] lut_15_table = 64'b0111011100000110011101010111011101000100000000000101010001110111;
    wire [5:0] lut_15_select = {
                             in_data[40],
                             in_data[39],
                             in_data[14],
                             in_data[30],
                             in_data[18],
                             in_data[38]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [63:0] lut_16_table = 64'b1100010000000000111111010000010011111100000000001111111100000100;
    wire [5:0] lut_16_select = {
                             in_data[56],
                             in_data[12],
                             in_data[52],
                             in_data[47],
                             in_data[46],
                             in_data[33]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [63:0] lut_17_table = 64'b0000000001000101111111111111111100000000010101010101111101111111;
    wire [5:0] lut_17_select = {
                             in_data[8],
                             in_data[17],
                             in_data[41],
                             in_data[49],
                             in_data[23],
                             in_data[13]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [63:0] lut_18_table = 64'b0000001001000010111111111101111101010011110111111111111111111111;
    wire [5:0] lut_18_select = {
                             in_data[42],
                             in_data[34],
                             in_data[54],
                             in_data[44],
                             in_data[29],
                             in_data[4]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [63:0] lut_19_table = 64'b1111001011111010111100001111101000100000111110100000000011111010;
    wire [5:0] lut_19_select = {
                             in_data[19],
                             in_data[48],
                             in_data[63],
                             in_data[31],
                             in_data[57],
                             in_data[0]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [63:0] lut_20_table = 64'b0011001100111011000100010011011100110111001010110001011100110111;
    wire [5:0] lut_20_select = {
                             in_data[60],
                             in_data[17],
                             in_data[62],
                             in_data[15],
                             in_data[7],
                             in_data[53]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [63:0] lut_21_table = 64'b1010111100101010001011110000101110001110000000000000111100001111;
    wire [5:0] lut_21_select = {
                             in_data[47],
                             in_data[0],
                             in_data[25],
                             in_data[5],
                             in_data[9],
                             in_data[63]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [63:0] lut_22_table = 64'b1111010111111111010100001101010101110001011101110101000001110101;
    wire [5:0] lut_22_select = {
                             in_data[43],
                             in_data[27],
                             in_data[45],
                             in_data[36],
                             in_data[51],
                             in_data[40]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [63:0] lut_23_table = 64'b1000110000001000100011110000101010001111100011111010111110101111;
    wire [5:0] lut_23_select = {
                             in_data[56],
                             in_data[18],
                             in_data[16],
                             in_data[6],
                             in_data[42],
                             in_data[21]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [63:0] lut_24_table = 64'b0011001110111111000000110000000000110011011101110011001100010011;
    wire [5:0] lut_24_select = {
                             in_data[41],
                             in_data[46],
                             in_data[57],
                             in_data[23],
                             in_data[49],
                             in_data[30]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [63:0] lut_25_table = 64'b0111000101010111111101011101010101010101010000010111010101010000;
    wire [5:0] lut_25_select = {
                             in_data[50],
                             in_data[52],
                             in_data[13],
                             in_data[12],
                             in_data[29],
                             in_data[59]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [63:0] lut_26_table = 64'b0101000101010101000001010000010101010101010111010001010000001101;
    wire [5:0] lut_26_select = {
                             in_data[33],
                             in_data[10],
                             in_data[54],
                             in_data[4],
                             in_data[48],
                             in_data[55]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [63:0] lut_27_table = 64'b0000110000001000110011001100110001001100010011000100110001000100;
    wire [5:0] lut_27_select = {
                             in_data[1],
                             in_data[37],
                             in_data[39],
                             in_data[26],
                             in_data[2],
                             in_data[58]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [63:0] lut_28_table = 64'b0111001111110111000000011101000100010001111101110000000101010001;
    wire [5:0] lut_28_select = {
                             in_data[11],
                             in_data[22],
                             in_data[32],
                             in_data[38],
                             in_data[34],
                             in_data[35]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [63:0] lut_29_table = 64'b1111110011111000111111111111110101001100000000000111011101110001;
    wire [5:0] lut_29_select = {
                             in_data[44],
                             in_data[61],
                             in_data[31],
                             in_data[8],
                             in_data[14],
                             in_data[3]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [63:0] lut_30_table = 64'b1111001111110111011101110011001100111111001101110000111100100011;
    wire [5:0] lut_30_select = {
                             in_data[57],
                             in_data[5],
                             in_data[20],
                             in_data[28],
                             in_data[19],
                             in_data[24]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [63:0] lut_31_table = 64'b1110111011111111110001001111111101001100010011000100010001000101;
    wire [5:0] lut_31_select = {
                             in_data[44],
                             in_data[38],
                             in_data[46],
                             in_data[18],
                             in_data[9],
                             in_data[61]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [63:0] lut_32_table = 64'b1111011111110000111101110110000001010101010001110111010100000000;
    wire [5:0] lut_32_select = {
                             in_data[21],
                             in_data[37],
                             in_data[29],
                             in_data[52],
                             in_data[60],
                             in_data[16]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [63:0] lut_33_table = 64'b0000000000000001000000000001011111111111010101111111111101111111;
    wire [5:0] lut_33_select = {
                             in_data[58],
                             in_data[54],
                             in_data[50],
                             in_data[35],
                             in_data[30],
                             in_data[4]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [63:0] lut_34_table = 64'b1110111111111111101011111111111111111111010101011110111111011111;
    wire [5:0] lut_34_select = {
                             in_data[34],
                             in_data[56],
                             in_data[31],
                             in_data[27],
                             in_data[43],
                             in_data[6]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [63:0] lut_35_table = 64'b0101111101011110111111101100110011111111111111101111111011111000;
    wire [5:0] lut_35_select = {
                             in_data[45],
                             in_data[0],
                             in_data[2],
                             in_data[3],
                             in_data[40],
                             in_data[15]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [63:0] lut_36_table = 64'b0111111111111111000100000011001000110111001100010000000000000000;
    wire [5:0] lut_36_select = {
                             in_data[26],
                             in_data[51],
                             in_data[22],
                             in_data[23],
                             in_data[49],
                             in_data[39]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [63:0] lut_37_table = 64'b1101100011111111100100000010100111111000111111111101100011111111;
    wire [5:0] lut_37_select = {
                             in_data[59],
                             in_data[55],
                             in_data[42],
                             in_data[48],
                             in_data[17],
                             in_data[36]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [63:0] lut_38_table = 64'b0010000011110001000100000111010100110000001100000001000001110001;
    wire [5:0] lut_38_select = {
                             in_data[41],
                             in_data[63],
                             in_data[10],
                             in_data[1],
                             in_data[7],
                             in_data[11]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [63:0] lut_39_table = 64'b0111011101110101011100110111010100010001010101010111001101110110;
    wire [5:0] lut_39_select = {
                             in_data[32],
                             in_data[62],
                             in_data[53],
                             in_data[8],
                             in_data[33],
                             in_data[25]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [63:0] lut_40_table = 64'b1111111110111111111110101010101010111110101011011010100010101000;
    wire [5:0] lut_40_select = {
                             in_data[0],
                             in_data[62],
                             in_data[14],
                             in_data[13],
                             in_data[47],
                             in_data[12]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [63:0] lut_41_table = 64'b0000000000000100000001001111110110001100100011001010100010111100;
    wire [5:0] lut_41_select = {
                             in_data[28],
                             in_data[9],
                             in_data[25],
                             in_data[50],
                             in_data[43],
                             in_data[37]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [63:0] lut_42_table = 64'b0010000000110000001100000011000010101010001000000111010000100000;
    wire [5:0] lut_42_select = {
                             in_data[61],
                             in_data[24],
                             in_data[29],
                             in_data[63],
                             in_data[56],
                             in_data[4]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [63:0] lut_43_table = 64'b0000100000001101000011000000110000011000000111011000110110001101;
    wire [5:0] lut_43_select = {
                             in_data[26],
                             in_data[30],
                             in_data[58],
                             in_data[49],
                             in_data[44],
                             in_data[53]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [63:0] lut_44_table = 64'b1011111100100011001011110000011110101111100000000000011100000000;
    wire [5:0] lut_44_select = {
                             in_data[34],
                             in_data[57],
                             in_data[16],
                             in_data[32],
                             in_data[20],
                             in_data[59]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [63:0] lut_45_table = 64'b0000010111011111000001011111111110001100101011110000100010101110;
    wire [5:0] lut_45_select = {
                             in_data[31],
                             in_data[23],
                             in_data[5],
                             in_data[18],
                             in_data[36],
                             in_data[51]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [63:0] lut_46_table = 64'b1010111011011101000000000000000011111110111111111010000011000000;
    wire [5:0] lut_46_select = {
                             in_data[46],
                             in_data[17],
                             in_data[11],
                             in_data[8],
                             in_data[1],
                             in_data[22]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [63:0] lut_47_table = 64'b1010011111111111100011001100111000110111111101111100111100000111;
    wire [5:0] lut_47_select = {
                             in_data[6],
                             in_data[21],
                             in_data[2],
                             in_data[45],
                             in_data[54],
                             in_data[60]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [63:0] lut_48_table = 64'b0000101000000000111111111111111000000000000000001110101011001000;
    wire [5:0] lut_48_select = {
                             in_data[39],
                             in_data[33],
                             in_data[41],
                             in_data[35],
                             in_data[10],
                             in_data[48]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [63:0] lut_49_table = 64'b0000000010101011000011110010111100000011001000110010101100101111;
    wire [5:0] lut_49_select = {
                             in_data[55],
                             in_data[15],
                             in_data[40],
                             in_data[42],
                             in_data[3],
                             in_data[52]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [63:0] lut_50_table = 64'b1110111011111010111010101111101011001000111110101100100011111010;
    wire [5:0] lut_50_select = {
                             in_data[46],
                             in_data[4],
                             in_data[19],
                             in_data[7],
                             in_data[27],
                             in_data[38]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [63:0] lut_51_table = 64'b1101110111001100110111001000100011011100000010001111110000000000;
    wire [5:0] lut_51_select = {
                             in_data[3],
                             in_data[47],
                             in_data[10],
                             in_data[23],
                             in_data[2],
                             in_data[51]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [63:0] lut_52_table = 64'b1011111111111111001111011111111100111101101111110001110111111111;
    wire [5:0] lut_52_select = {
                             in_data[12],
                             in_data[48],
                             in_data[57],
                             in_data[39],
                             in_data[44],
                             in_data[22]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [63:0] lut_53_table = 64'b0000101100001010100010111111111100000000000001000000000011111101;
    wire [5:0] lut_53_select = {
                             in_data[63],
                             in_data[34],
                             in_data[42],
                             in_data[40],
                             in_data[9],
                             in_data[54]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [63:0] lut_54_table = 64'b1100111100001000010111110000000011101111100011101110111100001000;
    wire [5:0] lut_54_select = {
                             in_data[16],
                             in_data[30],
                             in_data[18],
                             in_data[55],
                             in_data[60],
                             in_data[20]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [63:0] lut_55_table = 64'b1111101111111011000000001000000010001010101000001000000010100000;
    wire [5:0] lut_55_select = {
                             in_data[31],
                             in_data[26],
                             in_data[21],
                             in_data[62],
                             in_data[14],
                             in_data[56]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [63:0] lut_56_table = 64'b0010001000000010000000100000001011111010111111111111111111111111;
    wire [5:0] lut_56_select = {
                             in_data[61],
                             in_data[15],
                             in_data[8],
                             in_data[28],
                             in_data[32],
                             in_data[24]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [63:0] lut_57_table = 64'b0111011101110101111111111111011100110000111101010000000011010000;
    wire [5:0] lut_57_select = {
                             in_data[13],
                             in_data[11],
                             in_data[17],
                             in_data[5],
                             in_data[35],
                             in_data[43]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [63:0] lut_58_table = 64'b0000110011000000000000000000000001010101111111110000000001010000;
    wire [5:0] lut_58_select = {
                             in_data[41],
                             in_data[37],
                             in_data[53],
                             in_data[52],
                             in_data[33],
                             in_data[58]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [63:0] lut_59_table = 64'b0011111100001111011111110000111100001111000000100010111100000010;
    wire [5:0] lut_59_select = {
                             in_data[45],
                             in_data[50],
                             in_data[49],
                             in_data[6],
                             in_data[1],
                             in_data[29]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [63:0] lut_60_table = 64'b1111010111010101111111110000000011111111010101011111111100000100;
    wire [5:0] lut_60_select = {
                             in_data[63],
                             in_data[6],
                             in_data[25],
                             in_data[36],
                             in_data[0],
                             in_data[59]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [63:0] lut_61_table = 64'b0011001000110011101111110011111100110011000100110011111100011111;
    wire [5:0] lut_61_select = {
                             in_data[50],
                             in_data[30],
                             in_data[52],
                             in_data[53],
                             in_data[47],
                             in_data[20]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [63:0] lut_62_table = 64'b0000110011001101000001001100110011111111111111111111111111101110;
    wire [5:0] lut_62_select = {
                             in_data[35],
                             in_data[31],
                             in_data[48],
                             in_data[19],
                             in_data[4],
                             in_data[23]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [63:0] lut_63_table = 64'b0000111100001111101011101010111000001111000011110111101111101110;
    wire [5:0] lut_63_select = {
                             in_data[58],
                             in_data[28],
                             in_data[16],
                             in_data[62],
                             in_data[34],
                             in_data[26]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [63:0] lut_64_table = 64'b1111111011100000111110101110000011111010101000001110000011000000;
    wire [5:0] lut_64_select = {
                             in_data[42],
                             in_data[37],
                             in_data[15],
                             in_data[41],
                             in_data[5],
                             in_data[40]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [63:0] lut_65_table = 64'b0000000100000000110110010000000010111111000011111111111100001111;
    wire [5:0] lut_65_select = {
                             in_data[46],
                             in_data[21],
                             in_data[49],
                             in_data[12],
                             in_data[29],
                             in_data[44]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [63:0] lut_66_table = 64'b0101010100000101001101110000011101001111000000110000001100000011;
    wire [5:0] lut_66_select = {
                             in_data[32],
                             in_data[38],
                             in_data[55],
                             in_data[22],
                             in_data[51],
                             in_data[8]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [63:0] lut_67_table = 64'b1010101110001010111011111010101010001011100010101110111110101011;
    wire [5:0] lut_67_select = {
                             in_data[33],
                             in_data[39],
                             in_data[61],
                             in_data[2],
                             in_data[9],
                             in_data[54]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [63:0] lut_68_table = 64'b0010001100110011001000110011001100010011011100110101001101110011;
    wire [5:0] lut_68_select = {
                             in_data[3],
                             in_data[13],
                             in_data[7],
                             in_data[1],
                             in_data[24],
                             in_data[10]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [63:0] lut_69_table = 64'b0101000000010000011100010101000100010000000100000111001101110001;
    wire [5:0] lut_69_select = {
                             in_data[11],
                             in_data[45],
                             in_data[60],
                             in_data[43],
                             in_data[56],
                             in_data[18]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [63:0] lut_70_table = 64'b0000010000000000111111110001110100000000000000000011111100000000;
    wire [5:0] lut_70_select = {
                             in_data[35],
                             in_data[3],
                             in_data[57],
                             in_data[14],
                             in_data[27],
                             in_data[17]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [63:0] lut_71_table = 64'b0011111100111011111111111011011100101011001000100011101100110010;
    wire [5:0] lut_71_select = {
                             in_data[39],
                             in_data[62],
                             in_data[43],
                             in_data[28],
                             in_data[15],
                             in_data[41]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [63:0] lut_72_table = 64'b0100000011111111010000001111111100000000111000000000000011101110;
    wire [5:0] lut_72_select = {
                             in_data[53],
                             in_data[34],
                             in_data[32],
                             in_data[38],
                             in_data[33],
                             in_data[16]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [63:0] lut_73_table = 64'b1110111110101110111111111110111010101110100010001010100010001000;
    wire [5:0] lut_73_select = {
                             in_data[9],
                             in_data[61],
                             in_data[44],
                             in_data[12],
                             in_data[59],
                             in_data[6]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [63:0] lut_74_table = 64'b0000000000000000110111001101000011010100111100011111111111110111;
    wire [5:0] lut_74_select = {
                             in_data[18],
                             in_data[48],
                             in_data[7],
                             in_data[21],
                             in_data[8],
                             in_data[22]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [63:0] lut_75_table = 64'b1011111100000010001111110000001100111111000000100011111100000010;
    wire [5:0] lut_75_select = {
                             in_data[0],
                             in_data[11],
                             in_data[54],
                             in_data[5],
                             in_data[45],
                             in_data[29]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [63:0] lut_76_table = 64'b1010110001001100111111111111111100000000000000000010000001010000;
    wire [5:0] lut_76_select = {
                             in_data[23],
                             in_data[40],
                             in_data[46],
                             in_data[26],
                             in_data[25],
                             in_data[37]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [63:0] lut_77_table = 64'b0000101001011100000010001101110000001010000011000000110001001100;
    wire [5:0] lut_77_select = {
                             in_data[52],
                             in_data[24],
                             in_data[19],
                             in_data[31],
                             in_data[49],
                             in_data[56]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [63:0] lut_78_table = 64'b1011111100100010001110110010001011111111001010101011101100100010;
    wire [5:0] lut_78_select = {
                             in_data[50],
                             in_data[60],
                             in_data[4],
                             in_data[63],
                             in_data[30],
                             in_data[2]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [63:0] lut_79_table = 64'b0011001101110111000000010011000100111111011111110011001100110101;
    wire [5:0] lut_79_select = {
                             in_data[13],
                             in_data[58],
                             in_data[42],
                             in_data[55],
                             in_data[36],
                             in_data[47]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [63:0] lut_80_table = 64'b0000101000001000101110111011101110001011000010101111111110011111;
    wire [5:0] lut_80_select = {
                             in_data[6],
                             in_data[0],
                             in_data[1],
                             in_data[51],
                             in_data[20],
                             in_data[10]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [63:0] lut_81_table = 64'b1111101011111010111110100000001010000000000000001110100000000000;
    wire [5:0] lut_81_select = {
                             in_data[30],
                             in_data[12],
                             in_data[15],
                             in_data[26],
                             in_data[62],
                             in_data[48]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [63:0] lut_82_table = 64'b0101111100011011111111110111111101001111010111111100111111011111;
    wire [5:0] lut_82_select = {
                             in_data[19],
                             in_data[14],
                             in_data[4],
                             in_data[50],
                             in_data[53],
                             in_data[42]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [63:0] lut_83_table = 64'b0010001000000000001000100010001010101010111010001011101100100000;
    wire [5:0] lut_83_select = {
                             in_data[8],
                             in_data[32],
                             in_data[2],
                             in_data[33],
                             in_data[22],
                             in_data[31]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [63:0] lut_84_table = 64'b0000010100000101000011110001010100001111110011110000111110111111;
    wire [5:0] lut_84_select = {
                             in_data[39],
                             in_data[38],
                             in_data[35],
                             in_data[23],
                             in_data[7],
                             in_data[16]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [63:0] lut_85_table = 64'b0001000011010011000100011101111101110000100100001101001111111011;
    wire [5:0] lut_85_select = {
                             in_data[29],
                             in_data[43],
                             in_data[55],
                             in_data[63],
                             in_data[46],
                             in_data[5]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [63:0] lut_86_table = 64'b0100010011000100111111111110110100000000000000001111111111001101;
    wire [5:0] lut_86_select = {
                             in_data[24],
                             in_data[11],
                             in_data[41],
                             in_data[37],
                             in_data[21],
                             in_data[18]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [63:0] lut_87_table = 64'b0000111100001110000010000000100000001111100011110000111110101111;
    wire [5:0] lut_87_select = {
                             in_data[60],
                             in_data[54],
                             in_data[9],
                             in_data[45],
                             in_data[34],
                             in_data[58]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [63:0] lut_88_table = 64'b0000001100000000101010111010101001010001000000000111001100000010;
    wire [5:0] lut_88_select = {
                             in_data[56],
                             in_data[25],
                             in_data[27],
                             in_data[52],
                             in_data[49],
                             in_data[3]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [63:0] lut_89_table = 64'b1111000011111111110100001111111100000000111110110000000011000000;
    wire [5:0] lut_89_select = {
                             in_data[44],
                             in_data[47],
                             in_data[57],
                             in_data[59],
                             in_data[28],
                             in_data[17]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [63:0] lut_90_table = 64'b1100000001000010111000001010001000000000001010100000000000000010;
    wire [5:0] lut_90_select = {
                             in_data[57],
                             in_data[45],
                             in_data[36],
                             in_data[61],
                             in_data[13],
                             in_data[40]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [63:0] lut_91_table = 64'b1011000011111000100000001010100011111101111010001010101010101000;
    wire [5:0] lut_91_select = {
                             in_data[47],
                             in_data[4],
                             in_data[0],
                             in_data[30],
                             in_data[22],
                             in_data[49]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [63:0] lut_92_table = 64'b1100110011010101110011001100010011001100111111001100100011011100;
    wire [5:0] lut_92_select = {
                             in_data[10],
                             in_data[27],
                             in_data[29],
                             in_data[63],
                             in_data[59],
                             in_data[31]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [63:0] lut_93_table = 64'b1010111101100111111011101111111100000000000000000000000000000000;
    wire [5:0] lut_93_select = {
                             in_data[2],
                             in_data[15],
                             in_data[16],
                             in_data[44],
                             in_data[12],
                             in_data[50]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [63:0] lut_94_table = 64'b0011011110110011000000001011101000000000000000000000000000000000;
    wire [5:0] lut_94_select = {
                             in_data[32],
                             in_data[20],
                             in_data[17],
                             in_data[53],
                             in_data[51],
                             in_data[21]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [63:0] lut_95_table = 64'b1100111111011111111011111100111100001000000011001100111001001110;
    wire [5:0] lut_95_select = {
                             in_data[52],
                             in_data[58],
                             in_data[46],
                             in_data[37],
                             in_data[28],
                             in_data[26]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [63:0] lut_96_table = 64'b0011111100000011001110110011000000001011000000110000001000000000;
    wire [5:0] lut_96_select = {
                             in_data[62],
                             in_data[56],
                             in_data[55],
                             in_data[11],
                             in_data[8],
                             in_data[23]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [63:0] lut_97_table = 64'b1100111011101111101010101011101111001100100010111000000010111001;
    wire [5:0] lut_97_select = {
                             in_data[7],
                             in_data[3],
                             in_data[18],
                             in_data[38],
                             in_data[43],
                             in_data[6]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [63:0] lut_98_table = 64'b1010101010101111001000101010101010001010101011110000001010101010;
    wire [5:0] lut_98_select = {
                             in_data[24],
                             in_data[25],
                             in_data[14],
                             in_data[41],
                             in_data[39],
                             in_data[9]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [63:0] lut_99_table = 64'b1111111111110111001000100011001100000010000000000010101100111011;
    wire [5:0] lut_99_select = {
                             in_data[33],
                             in_data[35],
                             in_data[60],
                             in_data[19],
                             in_data[34],
                             in_data[1]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [63:0] lut_100_table = 64'b0000000011110111110101011111110100000000010101010100000001000100;
    wire [5:0] lut_100_select = {
                             in_data[57],
                             in_data[27],
                             in_data[54],
                             in_data[48],
                             in_data[5],
                             in_data[42]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [63:0] lut_101_table = 64'b1111111100101011101010100000000011111111101000101010001010100000;
    wire [5:0] lut_101_select = {
                             in_data[43],
                             in_data[10],
                             in_data[21],
                             in_data[25],
                             in_data[63],
                             in_data[22]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [63:0] lut_102_table = 64'b1110100011101000111010101111101010100000101000001110101011100000;
    wire [5:0] lut_102_select = {
                             in_data[11],
                             in_data[59],
                             in_data[35],
                             in_data[28],
                             in_data[38],
                             in_data[52]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [63:0] lut_103_table = 64'b1111001011110000111110101111111011100010110000001111101011111010;
    wire [5:0] lut_103_select = {
                             in_data[15],
                             in_data[19],
                             in_data[58],
                             in_data[9],
                             in_data[8],
                             in_data[61]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [63:0] lut_104_table = 64'b1000100010001000110011001111111110001000110011001100110011111111;
    wire [5:0] lut_104_select = {
                             in_data[17],
                             in_data[3],
                             in_data[33],
                             in_data[49],
                             in_data[62],
                             in_data[29]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [63:0] lut_105_table = 64'b0000000010000000101000001111100010001000101110111011101011111011;
    wire [5:0] lut_105_select = {
                             in_data[4],
                             in_data[51],
                             in_data[0],
                             in_data[39],
                             in_data[40],
                             in_data[34]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [63:0] lut_106_table = 64'b1110111010100010100011001010000010101110101010000000110000000100;
    wire [5:0] lut_106_select = {
                             in_data[23],
                             in_data[56],
                             in_data[1],
                             in_data[7],
                             in_data[37],
                             in_data[44]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [63:0] lut_107_table = 64'b1110101111111111000011101100111100001010100010100000001000000010;
    wire [5:0] lut_107_select = {
                             in_data[18],
                             in_data[12],
                             in_data[16],
                             in_data[53],
                             in_data[45],
                             in_data[60]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [63:0] lut_108_table = 64'b0000000001111101001100111111111100000000000001000011001011111111;
    wire [5:0] lut_108_select = {
                             in_data[13],
                             in_data[55],
                             in_data[14],
                             in_data[41],
                             in_data[47],
                             in_data[30]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [63:0] lut_109_table = 64'b0000101000001010101111111010111000000010000010100010101110101110;
    wire [5:0] lut_109_select = {
                             in_data[20],
                             in_data[26],
                             in_data[24],
                             in_data[50],
                             in_data[2],
                             in_data[6]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [63:0] lut_110_table = 64'b0100010001001100110111011101111100000100000001001101110101001101;
    wire [5:0] lut_110_select = {
                             in_data[48],
                             in_data[0],
                             in_data[46],
                             in_data[31],
                             in_data[32],
                             in_data[36]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [63:0] lut_111_table = 64'b1100000000000001110001000000000111000100000000001111110000000000;
    wire [5:0] lut_111_select = {
                             in_data[11],
                             in_data[53],
                             in_data[2],
                             in_data[58],
                             in_data[49],
                             in_data[39]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [63:0] lut_112_table = 64'b1101111111111111110001001101110111001100111111000100000011000100;
    wire [5:0] lut_112_select = {
                             in_data[9],
                             in_data[6],
                             in_data[13],
                             in_data[60],
                             in_data[59],
                             in_data[10]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [63:0] lut_113_table = 64'b0101111111011111000111110001000100011111010111010000000100000000;
    wire [5:0] lut_113_select = {
                             in_data[15],
                             in_data[17],
                             in_data[4],
                             in_data[43],
                             in_data[37],
                             in_data[25]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [63:0] lut_114_table = 64'b1110111100100010101011111011001011101111001000001011101100110000;
    wire [5:0] lut_114_select = {
                             in_data[38],
                             in_data[7],
                             in_data[29],
                             in_data[27],
                             in_data[47],
                             in_data[18]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [63:0] lut_115_table = 64'b1010111011111111000010001000111000111011111111110000000010001111;
    wire [5:0] lut_115_select = {
                             in_data[33],
                             in_data[14],
                             in_data[54],
                             in_data[8],
                             in_data[5],
                             in_data[1]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [63:0] lut_116_table = 64'b0111010100100000100011111010111100010001001000110000000000000010;
    wire [5:0] lut_116_select = {
                             in_data[50],
                             in_data[19],
                             in_data[24],
                             in_data[44],
                             in_data[3],
                             in_data[12]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [63:0] lut_117_table = 64'b1111011101010101111111110000010101110001000000011111011100000001;
    wire [5:0] lut_117_select = {
                             in_data[28],
                             in_data[57],
                             in_data[61],
                             in_data[35],
                             in_data[45],
                             in_data[63]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [63:0] lut_118_table = 64'b0000000000000000001000100010000000101010000010001011111111111111;
    wire [5:0] lut_118_select = {
                             in_data[52],
                             in_data[55],
                             in_data[56],
                             in_data[16],
                             in_data[62],
                             in_data[40]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [63:0] lut_119_table = 64'b0000000001010100000000001111110100000000011101000101000011111101;
    wire [5:0] lut_119_select = {
                             in_data[21],
                             in_data[34],
                             in_data[26],
                             in_data[30],
                             in_data[20],
                             in_data[23]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [63:0] lut_120_table = 64'b0100010111011101010011111100111101010101110101011100111111001101;
    wire [5:0] lut_120_select = {
                             in_data[29],
                             in_data[15],
                             in_data[51],
                             in_data[22],
                             in_data[41],
                             in_data[42]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [63:0] lut_121_table = 64'b0011001101110011001100110011001100000000000100110001000100010011;
    wire [5:0] lut_121_select = {
                             in_data[43],
                             in_data[48],
                             in_data[58],
                             in_data[39],
                             in_data[31],
                             in_data[21]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [63:0] lut_122_table = 64'b0100011111001111010001001100111101010011110101111101011111111111;
    wire [5:0] lut_122_select = {
                             in_data[37],
                             in_data[28],
                             in_data[16],
                             in_data[27],
                             in_data[53],
                             in_data[8]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [63:0] lut_123_table = 64'b1101110000000000110011110000100011011110000010001110111100101010;
    wire [5:0] lut_123_select = {
                             in_data[14],
                             in_data[56],
                             in_data[10],
                             in_data[46],
                             in_data[60],
                             in_data[3]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [63:0] lut_124_table = 64'b0011001001110011011100001111000011111111111111111111001011111111;
    wire [5:0] lut_124_select = {
                             in_data[17],
                             in_data[23],
                             in_data[33],
                             in_data[19],
                             in_data[1],
                             in_data[6]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [63:0] lut_125_table = 64'b1100110111111111110111111111111111011111111110111101111111110010;
    wire [5:0] lut_125_select = {
                             in_data[34],
                             in_data[38],
                             in_data[55],
                             in_data[36],
                             in_data[59],
                             in_data[7]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [63:0] lut_126_table = 64'b0000000001011111000000000100111100000010111111110000011001111111;
    wire [5:0] lut_126_select = {
                             in_data[35],
                             in_data[49],
                             in_data[25],
                             in_data[57],
                             in_data[24],
                             in_data[20]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [63:0] lut_127_table = 64'b1111011111111111111100001000100000110011000000110111000000000000;
    wire [5:0] lut_127_select = {
                             in_data[9],
                             in_data[32],
                             in_data[11],
                             in_data[40],
                             in_data[62],
                             in_data[45]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [63:0] lut_128_table = 64'b0000000100000011001000110010001111001111100011111111111110101111;
    wire [5:0] lut_128_select = {
                             in_data[52],
                             in_data[50],
                             in_data[0],
                             in_data[12],
                             in_data[63],
                             in_data[2]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [63:0] lut_129_table = 64'b1111111111111111000010001111101101001111010111110000100000001010;
    wire [5:0] lut_129_select = {
                             in_data[54],
                             in_data[26],
                             in_data[61],
                             in_data[44],
                             in_data[30],
                             in_data[47]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [63:0] lut_130_table = 64'b1010111100101111101010110010101010111111001011110011101000100011;
    wire [5:0] lut_130_select = {
                             in_data[41],
                             in_data[2],
                             in_data[13],
                             in_data[18],
                             in_data[5],
                             in_data[4]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [63:0] lut_131_table = 64'b1011111100110011101110111011001100000011000000100011001100000011;
    wire [5:0] lut_131_select = {
                             in_data[24],
                             in_data[30],
                             in_data[44],
                             in_data[39],
                             in_data[20],
                             in_data[59]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [63:0] lut_132_table = 64'b0000000000011011000001000011101100010000000111111111111111111111;
    wire [5:0] lut_132_select = {
                             in_data[3],
                             in_data[27],
                             in_data[55],
                             in_data[33],
                             in_data[38],
                             in_data[10]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [63:0] lut_133_table = 64'b0011000000010000000000001111101000001000000010001000101011111010;
    wire [5:0] lut_133_select = {
                             in_data[15],
                             in_data[19],
                             in_data[6],
                             in_data[51],
                             in_data[12],
                             in_data[57]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [63:0] lut_134_table = 64'b1111000011111010111111110100111011111100110111101111111100001100;
    wire [5:0] lut_134_select = {
                             in_data[54],
                             in_data[31],
                             in_data[50],
                             in_data[43],
                             in_data[63],
                             in_data[37]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [63:0] lut_135_table = 64'b1000110000000000111111111111110000000100000000001111110111111110;
    wire [5:0] lut_135_select = {
                             in_data[40],
                             in_data[61],
                             in_data[35],
                             in_data[52],
                             in_data[21],
                             in_data[28]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [63:0] lut_136_table = 64'b0111011101000000111111111111111000110011010000000111011101111110;
    wire [5:0] lut_136_select = {
                             in_data[32],
                             in_data[8],
                             in_data[34],
                             in_data[36],
                             in_data[16],
                             in_data[7]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [63:0] lut_137_table = 64'b0000101110101010000000100000000011111111111111110000011100100011;
    wire [5:0] lut_137_select = {
                             in_data[42],
                             in_data[45],
                             in_data[0],
                             in_data[62],
                             in_data[47],
                             in_data[58]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [63:0] lut_138_table = 64'b1100110001111111010011000101111111001100110111010100010011000100;
    wire [5:0] lut_138_select = {
                             in_data[22],
                             in_data[25],
                             in_data[14],
                             in_data[17],
                             in_data[60],
                             in_data[1]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [63:0] lut_139_table = 64'b0111001100000011001100110000001000110011000000100011001100000010;
    wire [5:0] lut_139_select = {
                             in_data[48],
                             in_data[23],
                             in_data[11],
                             in_data[9],
                             in_data[53],
                             in_data[29]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [63:0] lut_140_table = 64'b1111010011111100000000000000000011111110111111110001000001000101;
    wire [5:0] lut_140_select = {
                             in_data[48],
                             in_data[27],
                             in_data[46],
                             in_data[26],
                             in_data[49],
                             in_data[56]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [63:0] lut_141_table = 64'b1111110111111101110101010000010011010100010001000000010000000100;
    wire [5:0] lut_141_select = {
                             in_data[45],
                             in_data[3],
                             in_data[43],
                             in_data[35],
                             in_data[53],
                             in_data[0]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [63:0] lut_142_table = 64'b1011101100110010101100001011101011110001001100100011000001110000;
    wire [5:0] lut_142_select = {
                             in_data[17],
                             in_data[37],
                             in_data[58],
                             in_data[24],
                             in_data[47],
                             in_data[16]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [63:0] lut_143_table = 64'b0111010100000000010101000000010011110111011101010111010101110101;
    wire [5:0] lut_143_select = {
                             in_data[60],
                             in_data[2],
                             in_data[38],
                             in_data[59],
                             in_data[25],
                             in_data[62]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [63:0] lut_144_table = 64'b1011111100101111101100110010001100000010000000100000000000000000;
    wire [5:0] lut_144_select = {
                             in_data[19],
                             in_data[14],
                             in_data[13],
                             in_data[11],
                             in_data[52],
                             in_data[23]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [63:0] lut_145_table = 64'b1111011111110101110000001101000011110010111101010010000001000000;
    wire [5:0] lut_145_select = {
                             in_data[32],
                             in_data[8],
                             in_data[21],
                             in_data[20],
                             in_data[51],
                             in_data[30]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [63:0] lut_146_table = 64'b1100010000000100110000000000000011110100111111011100010011010100;
    wire [5:0] lut_146_select = {
                             in_data[4],
                             in_data[7],
                             in_data[18],
                             in_data[55],
                             in_data[28],
                             in_data[9]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [63:0] lut_147_table = 64'b1111111111001100111111111110110011001100110011001100110010001000;
    wire [5:0] lut_147_select = {
                             in_data[54],
                             in_data[50],
                             in_data[15],
                             in_data[33],
                             in_data[31],
                             in_data[40]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [63:0] lut_148_table = 64'b0000111000001100000010101000111011101110111011001000101011101110;
    wire [5:0] lut_148_select = {
                             in_data[63],
                             in_data[1],
                             in_data[34],
                             in_data[22],
                             in_data[36],
                             in_data[10]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [63:0] lut_149_table = 64'b0000101110001111000010111001101110111111111111111011111110111011;
    wire [5:0] lut_149_select = {
                             in_data[44],
                             in_data[39],
                             in_data[61],
                             in_data[57],
                             in_data[42],
                             in_data[5]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [63:0] lut_150_table = 64'b0000000000000000000000000100111110000000111010001010100011111111;
    wire [5:0] lut_150_select = {
                             in_data[31],
                             in_data[14],
                             in_data[29],
                             in_data[41],
                             in_data[12],
                             in_data[6]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [63:0] lut_151_table = 64'b0101000011110100000100001111010001010100111111110101010111111111;
    wire [5:0] lut_151_select = {
                             in_data[30],
                             in_data[46],
                             in_data[40],
                             in_data[38],
                             in_data[34],
                             in_data[3]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [63:0] lut_152_table = 64'b1111111111110000111111111111000011110111010100000111011101010000;
    wire [5:0] lut_152_select = {
                             in_data[1],
                             in_data[8],
                             in_data[5],
                             in_data[56],
                             in_data[43],
                             in_data[28]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [63:0] lut_153_table = 64'b1101000011111100000000000000000011111000111111000000000011010100;
    wire [5:0] lut_153_select = {
                             in_data[15],
                             in_data[62],
                             in_data[24],
                             in_data[32],
                             in_data[27],
                             in_data[50]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [63:0] lut_154_table = 64'b0000000000110011001000001011001000100010001100110010001010110011;
    wire [5:0] lut_154_select = {
                             in_data[18],
                             in_data[59],
                             in_data[58],
                             in_data[61],
                             in_data[21],
                             in_data[37]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [63:0] lut_155_table = 64'b0000000010101010000000101010111100000000111011100000001011101111;
    wire [5:0] lut_155_select = {
                             in_data[23],
                             in_data[39],
                             in_data[48],
                             in_data[44],
                             in_data[36],
                             in_data[42]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [63:0] lut_156_table = 64'b0000000001110101000000100011011100000000011101110011001101111111;
    wire [5:0] lut_156_select = {
                             in_data[63],
                             in_data[16],
                             in_data[9],
                             in_data[45],
                             in_data[57],
                             in_data[35]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [63:0] lut_157_table = 64'b1100111110001100111111111100111110001111000000001111111110001111;
    wire [5:0] lut_157_select = {
                             in_data[20],
                             in_data[47],
                             in_data[52],
                             in_data[53],
                             in_data[54],
                             in_data[2]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [63:0] lut_158_table = 64'b1111111101010000010100010000000011111111000100001111111100000000;
    wire [5:0] lut_158_select = {
                             in_data[19],
                             in_data[33],
                             in_data[60],
                             in_data[13],
                             in_data[26],
                             in_data[7]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [63:0] lut_159_table = 64'b1011111110001011101110110010001100000000000000000000000100110011;
    wire [5:0] lut_159_select = {
                             in_data[25],
                             in_data[4],
                             in_data[11],
                             in_data[49],
                             in_data[51],
                             in_data[22]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [63:0] lut_160_table = 64'b1111000011110010000000000101000011110000111110110101000011110000;
    wire [5:0] lut_160_select = {
                             in_data[30],
                             in_data[20],
                             in_data[10],
                             in_data[17],
                             in_data[55],
                             in_data[0]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [63:0] lut_161_table = 64'b0010101110111010001100001111111100000000000100000000000001010000;
    wire [5:0] lut_161_select = {
                             in_data[58],
                             in_data[57],
                             in_data[44],
                             in_data[50],
                             in_data[28],
                             in_data[61]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [63:0] lut_162_table = 64'b0000000101010101000000010101010110000101111111011000110111111101;
    wire [5:0] lut_162_select = {
                             in_data[36],
                             in_data[23],
                             in_data[32],
                             in_data[37],
                             in_data[48],
                             in_data[18]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [63:0] lut_163_table = 64'b1110110111101111111111111111111100000000000000000001000100000001;
    wire [5:0] lut_163_select = {
                             in_data[53],
                             in_data[49],
                             in_data[8],
                             in_data[5],
                             in_data[11],
                             in_data[38]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [63:0] lut_164_table = 64'b0101000001110000010100000101000011110101111101110111000101010001;
    wire [5:0] lut_164_select = {
                             in_data[35],
                             in_data[3],
                             in_data[59],
                             in_data[21],
                             in_data[33],
                             in_data[45]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [63:0] lut_165_table = 64'b1010001011101111111011111110111100100011111001111110111111101111;
    wire [5:0] lut_165_select = {
                             in_data[62],
                             in_data[16],
                             in_data[15],
                             in_data[54],
                             in_data[19],
                             in_data[39]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [63:0] lut_166_table = 64'b1011111110111111000000110000001111111111111111110000001100001111;
    wire [5:0] lut_166_select = {
                             in_data[2],
                             in_data[29],
                             in_data[7],
                             in_data[13],
                             in_data[51],
                             in_data[26]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [63:0] lut_167_table = 64'b1111111101110011011111110001001001011111000000000100111100000000;
    wire [5:0] lut_167_select = {
                             in_data[25],
                             in_data[43],
                             in_data[47],
                             in_data[42],
                             in_data[60],
                             in_data[6]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [63:0] lut_168_table = 64'b1100111110000000000000001000000011111111110011001100110011000000;
    wire [5:0] lut_168_select = {
                             in_data[40],
                             in_data[27],
                             in_data[22],
                             in_data[24],
                             in_data[1],
                             in_data[31]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [63:0] lut_169_table = 64'b1111101010101000110111001100010011101010101011101110111110001110;
    wire [5:0] lut_169_select = {
                             in_data[9],
                             in_data[4],
                             in_data[63],
                             in_data[41],
                             in_data[52],
                             in_data[12]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [63:0] lut_170_table = 64'b0010111110111111101010101010111110101111101011111000101010101011;
    wire [5:0] lut_170_select = {
                             in_data[17],
                             in_data[24],
                             in_data[46],
                             in_data[56],
                             in_data[14],
                             in_data[34]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [63:0] lut_171_table = 64'b0000000110110011000100111111111100000011000000010000101100110011;
    wire [5:0] lut_171_select = {
                             in_data[59],
                             in_data[4],
                             in_data[36],
                             in_data[40],
                             in_data[49],
                             in_data[5]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [63:0] lut_172_table = 64'b0011001110111011001000101111101100100010001010100000000000100010;
    wire [5:0] lut_172_select = {
                             in_data[12],
                             in_data[8],
                             in_data[23],
                             in_data[37],
                             in_data[0],
                             in_data[57]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [63:0] lut_173_table = 64'b1111111111111111111110101111111101010000010100000000000001110000;
    wire [5:0] lut_173_select = {
                             in_data[22],
                             in_data[10],
                             in_data[7],
                             in_data[16],
                             in_data[18],
                             in_data[42]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [63:0] lut_174_table = 64'b0000000011111111000000000000011100000000011001000100010001001101;
    wire [5:0] lut_174_select = {
                             in_data[19],
                             in_data[45],
                             in_data[52],
                             in_data[11],
                             in_data[6],
                             in_data[38]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [63:0] lut_175_table = 64'b0101010100000000111111111111111101010000000000000111010101010000;
    wire [5:0] lut_175_select = {
                             in_data[9],
                             in_data[33],
                             in_data[20],
                             in_data[15],
                             in_data[28],
                             in_data[27]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [63:0] lut_176_table = 64'b1010101010000010111011101000001010001010100010101100110011001110;
    wire [5:0] lut_176_select = {
                             in_data[53],
                             in_data[3],
                             in_data[55],
                             in_data[61],
                             in_data[35],
                             in_data[32]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [63:0] lut_177_table = 64'b1111110111011101110011001100010011001100110011000100000000000000;
    wire [5:0] lut_177_select = {
                             in_data[47],
                             in_data[25],
                             in_data[63],
                             in_data[39],
                             in_data[1],
                             in_data[60]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [63:0] lut_178_table = 64'b0000100011101100110010001000100011111111111111111110110010101000;
    wire [5:0] lut_178_select = {
                             in_data[54],
                             in_data[29],
                             in_data[31],
                             in_data[13],
                             in_data[62],
                             in_data[58]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [63:0] lut_179_table = 64'b0000000011111111000000001111111100000000111111110000001011111111;
    wire [5:0] lut_179_select = {
                             in_data[44],
                             in_data[21],
                             in_data[41],
                             in_data[26],
                             in_data[50],
                             in_data[48]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [63:0] lut_180_table = 64'b0100111100000100010011110000010011111111110011111111111101011111;
    wire [5:0] lut_180_select = {
                             in_data[34],
                             in_data[1],
                             in_data[43],
                             in_data[2],
                             in_data[30],
                             in_data[51]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [63:0] lut_181_table = 64'b1111110011011101110100001101110110000000100110000000000000010101;
    wire [5:0] lut_181_select = {
                             in_data[26],
                             in_data[5],
                             in_data[16],
                             in_data[45],
                             in_data[33],
                             in_data[57]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [63:0] lut_182_table = 64'b1111111110000000111111111111111100000000000000001111111111011101;
    wire [5:0] lut_182_select = {
                             in_data[44],
                             in_data[58],
                             in_data[8],
                             in_data[25],
                             in_data[10],
                             in_data[14]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [63:0] lut_183_table = 64'b1110111011101010101011101110111010100001001100001000110010100000;
    wire [5:0] lut_183_select = {
                             in_data[60],
                             in_data[41],
                             in_data[7],
                             in_data[62],
                             in_data[38],
                             in_data[31]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [63:0] lut_184_table = 64'b1111111101111111010011110100111100000111000011110000000000000000;
    wire [5:0] lut_184_select = {
                             in_data[3],
                             in_data[13],
                             in_data[4],
                             in_data[59],
                             in_data[56],
                             in_data[32]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [63:0] lut_185_table = 64'b1110111110001000111111111010000011101010101010001111101110101010;
    wire [5:0] lut_185_select = {
                             in_data[42],
                             in_data[22],
                             in_data[29],
                             in_data[11],
                             in_data[23],
                             in_data[28]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [63:0] lut_186_table = 64'b0011000000010000101010000000100000110000000100001011100000001000;
    wire [5:0] lut_186_select = {
                             in_data[54],
                             in_data[40],
                             in_data[24],
                             in_data[17],
                             in_data[36],
                             in_data[21]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [63:0] lut_187_table = 64'b0001100000110000100110100011001110011000111110100011100011110011;
    wire [5:0] lut_187_select = {
                             in_data[55],
                             in_data[37],
                             in_data[50],
                             in_data[39],
                             in_data[0],
                             in_data[19]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [63:0] lut_188_table = 64'b0100010111111111010001001111110000000100010001010000000011000100;
    wire [5:0] lut_188_select = {
                             in_data[61],
                             in_data[46],
                             in_data[20],
                             in_data[53],
                             in_data[48],
                             in_data[18]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [63:0] lut_189_table = 64'b0101111011111110111111111111111100000010000011100000001001001110;
    wire [5:0] lut_189_select = {
                             in_data[6],
                             in_data[35],
                             in_data[47],
                             in_data[12],
                             in_data[27],
                             in_data[63]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [63:0] lut_190_table = 64'b0101010100000000111111110100111101001100000010001111111111001111;
    wire [5:0] lut_190_select = {
                             in_data[17],
                             in_data[50],
                             in_data[9],
                             in_data[15],
                             in_data[49],
                             in_data[52]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [63:0] lut_191_table = 64'b0010000000000010111010101010101110100000001000001111101000111011;
    wire [5:0] lut_191_select = {
                             in_data[1],
                             in_data[4],
                             in_data[23],
                             in_data[27],
                             in_data[61],
                             in_data[32]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [63:0] lut_192_table = 64'b1111111011111100111111001100010011111100111011001100100011000000;
    wire [5:0] lut_192_select = {
                             in_data[58],
                             in_data[31],
                             in_data[55],
                             in_data[3],
                             in_data[0],
                             in_data[18]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [63:0] lut_193_table = 64'b0000010100001100010011111100011100000100100011000000010100000000;
    wire [5:0] lut_193_select = {
                             in_data[20],
                             in_data[60],
                             in_data[2],
                             in_data[7],
                             in_data[62],
                             in_data[36]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [63:0] lut_194_table = 64'b0000000011110101000000000101010001010001011101010101010111110101;
    wire [5:0] lut_194_select = {
                             in_data[43],
                             in_data[28],
                             in_data[57],
                             in_data[40],
                             in_data[26],
                             in_data[25]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [63:0] lut_195_table = 64'b0111010100000100010001010000010001011101010001010100110101000100;
    wire [5:0] lut_195_select = {
                             in_data[35],
                             in_data[24],
                             in_data[63],
                             in_data[13],
                             in_data[8],
                             in_data[19]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [63:0] lut_196_table = 64'b0001001100010011000010110011101100111111001111110011111100111111;
    wire [5:0] lut_196_select = {
                             in_data[34],
                             in_data[29],
                             in_data[56],
                             in_data[44],
                             in_data[53],
                             in_data[21]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [63:0] lut_197_table = 64'b0000000000010000000000001011000011011101111111110010010111111111;
    wire [5:0] lut_197_select = {
                             in_data[10],
                             in_data[59],
                             in_data[41],
                             in_data[51],
                             in_data[37],
                             in_data[38]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [63:0] lut_198_table = 64'b1011001010111010101100101011101010100010101100101011001010110010;
    wire [5:0] lut_198_select = {
                             in_data[33],
                             in_data[6],
                             in_data[16],
                             in_data[45],
                             in_data[22],
                             in_data[11]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [63:0] lut_199_table = 64'b1011111100110011101111110000000011111111000100011111111100000000;
    wire [5:0] lut_199_select = {
                             in_data[42],
                             in_data[5],
                             in_data[14],
                             in_data[47],
                             in_data[54],
                             in_data[48]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [63:0] lut_200_table = 64'b1111111111110000111111110111000011111111111100011111111111110111;
    wire [5:0] lut_200_select = {
                             in_data[23],
                             in_data[47],
                             in_data[30],
                             in_data[12],
                             in_data[39],
                             in_data[46]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [63:0] lut_201_table = 64'b1111111110101010111011111010001011111111101000101111111110111011;
    wire [5:0] lut_201_select = {
                             in_data[48],
                             in_data[51],
                             in_data[19],
                             in_data[3],
                             in_data[22],
                             in_data[44]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [63:0] lut_202_table = 64'b0000100000110011000011001011101000001000000000000000110000001000;
    wire [5:0] lut_202_select = {
                             in_data[11],
                             in_data[25],
                             in_data[2],
                             in_data[35],
                             in_data[14],
                             in_data[53]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [63:0] lut_203_table = 64'b0001000100010011000100000000000101111111101111110001000100110011;
    wire [5:0] lut_203_select = {
                             in_data[26],
                             in_data[1],
                             in_data[4],
                             in_data[29],
                             in_data[55],
                             in_data[31]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [63:0] lut_204_table = 64'b1110111010101110100011101110111100111110001011101110111111111111;
    wire [5:0] lut_204_select = {
                             in_data[27],
                             in_data[58],
                             in_data[16],
                             in_data[50],
                             in_data[56],
                             in_data[43]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [63:0] lut_205_table = 64'b0000001100000011000101110000000100000011000000110101011100010111;
    wire [5:0] lut_205_select = {
                             in_data[63],
                             in_data[62],
                             in_data[6],
                             in_data[52],
                             in_data[60],
                             in_data[13]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [63:0] lut_206_table = 64'b0000000001010101000000000001110100000000000111110000001101111111;
    wire [5:0] lut_206_select = {
                             in_data[34],
                             in_data[42],
                             in_data[5],
                             in_data[38],
                             in_data[37],
                             in_data[17]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [63:0] lut_207_table = 64'b1111110111111101110001001100010010110011111110111111000111110101;
    wire [5:0] lut_207_select = {
                             in_data[28],
                             in_data[59],
                             in_data[8],
                             in_data[32],
                             in_data[9],
                             in_data[7]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [63:0] lut_208_table = 64'b1111011100000001111101110111011111100100010000001100010001010101;
    wire [5:0] lut_208_select = {
                             in_data[24],
                             in_data[40],
                             in_data[20],
                             in_data[33],
                             in_data[10],
                             in_data[61]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [63:0] lut_209_table = 64'b1010111110001111000010100000111110001111100011110000101010001110;
    wire [5:0] lut_209_select = {
                             in_data[45],
                             in_data[36],
                             in_data[15],
                             in_data[41],
                             in_data[18],
                             in_data[0]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [63:0] lut_210_table = 64'b0010000000000000001100100101000010110000011100001111101111111101;
    wire [5:0] lut_210_select = {
                             in_data[11],
                             in_data[13],
                             in_data[21],
                             in_data[49],
                             in_data[57],
                             in_data[54]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [63:0] lut_211_table = 64'b1100110011001110110011001100100010001000111010101010100010101000;
    wire [5:0] lut_211_select = {
                             in_data[33],
                             in_data[12],
                             in_data[23],
                             in_data[59],
                             in_data[17],
                             in_data[6]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [63:0] lut_212_table = 64'b1111111111111111111100001111101000110000000100000010000010110000;
    wire [5:0] lut_212_select = {
                             in_data[3],
                             in_data[44],
                             in_data[52],
                             in_data[2],
                             in_data[61],
                             in_data[53]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [63:0] lut_213_table = 64'b1010001010100010101000101111101110100010101000101010000010111010;
    wire [5:0] lut_213_select = {
                             in_data[39],
                             in_data[14],
                             in_data[26],
                             in_data[20],
                             in_data[24],
                             in_data[63]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [63:0] lut_214_table = 64'b1111111110111111111111111011111100000011000001110000001100000111;
    wire [5:0] lut_214_select = {
                             in_data[60],
                             in_data[31],
                             in_data[25],
                             in_data[8],
                             in_data[19],
                             in_data[38]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [63:0] lut_215_table = 64'b1100010001000100111011101100111100000000010001001110100001000100;
    wire [5:0] lut_215_select = {
                             in_data[45],
                             in_data[10],
                             in_data[55],
                             in_data[58],
                             in_data[5],
                             in_data[28]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [63:0] lut_216_table = 64'b1111101100110010111100100010000011111011001000101011001000000000;
    wire [5:0] lut_216_select = {
                             in_data[29],
                             in_data[35],
                             in_data[42],
                             in_data[7],
                             in_data[43],
                             in_data[4]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [63:0] lut_217_table = 64'b1111111111111111111111011111111100000000111111110000000000000000;
    wire [5:0] lut_217_select = {
                             in_data[22],
                             in_data[9],
                             in_data[41],
                             in_data[1],
                             in_data[37],
                             in_data[15]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [63:0] lut_218_table = 64'b1010101010001000101011110000000011111010111100001111111111110111;
    wire [5:0] lut_218_select = {
                             in_data[0],
                             in_data[16],
                             in_data[56],
                             in_data[40],
                             in_data[48],
                             in_data[32]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [63:0] lut_219_table = 64'b0000000011101111000000000000101100001011111111110000101111111111;
    wire [5:0] lut_219_select = {
                             in_data[36],
                             in_data[51],
                             in_data[62],
                             in_data[47],
                             in_data[18],
                             in_data[34]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [63:0] lut_220_table = 64'b0100100011111111111011101111111100000000010100110000110000001100;
    wire [5:0] lut_220_select = {
                             in_data[59],
                             in_data[23],
                             in_data[50],
                             in_data[46],
                             in_data[27],
                             in_data[30]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [63:0] lut_221_table = 64'b1010101000100000100011100000000000001000101101000000101000000100;
    wire [5:0] lut_221_select = {
                             in_data[56],
                             in_data[29],
                             in_data[53],
                             in_data[26],
                             in_data[8],
                             in_data[21]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [63:0] lut_222_table = 64'b1000100010101010110011001110111011111010101010101100110010101110;
    wire [5:0] lut_222_select = {
                             in_data[9],
                             in_data[11],
                             in_data[51],
                             in_data[28],
                             in_data[39],
                             in_data[42]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [63:0] lut_223_table = 64'b0101111111111111000000010000000000100011111010110000000000000000;
    wire [5:0] lut_223_select = {
                             in_data[3],
                             in_data[2],
                             in_data[17],
                             in_data[47],
                             in_data[36],
                             in_data[63]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [63:0] lut_224_table = 64'b1111010001000100010011111111110001111111111101000000111100001110;
    wire [5:0] lut_224_select = {
                             in_data[62],
                             in_data[43],
                             in_data[60],
                             in_data[54],
                             in_data[57],
                             in_data[25]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [63:0] lut_225_table = 64'b1011000010110000101010100010000000000000101110100000100000001010;
    wire [5:0] lut_225_select = {
                             in_data[34],
                             in_data[45],
                             in_data[4],
                             in_data[35],
                             in_data[16],
                             in_data[32]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [63:0] lut_226_table = 64'b1010101010101010111110111111001100001010001010101010101011110011;
    wire [5:0] lut_226_select = {
                             in_data[48],
                             in_data[38],
                             in_data[18],
                             in_data[40],
                             in_data[37],
                             in_data[19]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [63:0] lut_227_table = 64'b1111001100110011000100110000001111111111111110111111001110110011;
    wire [5:0] lut_227_select = {
                             in_data[1],
                             in_data[49],
                             in_data[0],
                             in_data[33],
                             in_data[20],
                             in_data[52]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [63:0] lut_228_table = 64'b0000000000001100100011111100111100000110100011110000011111001111;
    wire [5:0] lut_228_select = {
                             in_data[5],
                             in_data[31],
                             in_data[55],
                             in_data[7],
                             in_data[58],
                             in_data[44]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [63:0] lut_229_table = 64'b0111001101110011010100000011000011111111111100111111001100110011;
    wire [5:0] lut_229_select = {
                             in_data[24],
                             in_data[61],
                             in_data[15],
                             in_data[13],
                             in_data[22],
                             in_data[10]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [63:0] lut_230_table = 64'b0000100000001111001110010011111100100000000010001011000000101011;
    wire [5:0] lut_230_select = {
                             in_data[25],
                             in_data[32],
                             in_data[41],
                             in_data[14],
                             in_data[12],
                             in_data[6]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [63:0] lut_231_table = 64'b1010001010110010000000000000000011111011111111111011001010110011;
    wire [5:0] lut_231_select = {
                             in_data[13],
                             in_data[0],
                             in_data[52],
                             in_data[49],
                             in_data[44],
                             in_data[19]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [63:0] lut_232_table = 64'b0000001100000000110000001100101000000001000000000000000010101011;
    wire [5:0] lut_232_select = {
                             in_data[57],
                             in_data[59],
                             in_data[9],
                             in_data[35],
                             in_data[21],
                             in_data[28]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [63:0] lut_233_table = 64'b0000000001010001110101001101010100001100010101011100110011011101;
    wire [5:0] lut_233_select = {
                             in_data[34],
                             in_data[63],
                             in_data[62],
                             in_data[42],
                             in_data[48],
                             in_data[50]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [63:0] lut_234_table = 64'b0000010100001101000000000100110111011111010101010000010100000101;
    wire [5:0] lut_234_select = {
                             in_data[18],
                             in_data[36],
                             in_data[7],
                             in_data[54],
                             in_data[8],
                             in_data[27]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [63:0] lut_235_table = 64'b1010100010110011110010111111111100100011001100110000001110111111;
    wire [5:0] lut_235_select = {
                             in_data[43],
                             in_data[10],
                             in_data[47],
                             in_data[33],
                             in_data[2],
                             in_data[39]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [63:0] lut_236_table = 64'b1111011111111111011100110011001100110011001100010001000100000000;
    wire [5:0] lut_236_select = {
                             in_data[31],
                             in_data[1],
                             in_data[5],
                             in_data[53],
                             in_data[22],
                             in_data[30]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [63:0] lut_237_table = 64'b0000000000000100000000001111010101111111011111111111111111111111;
    wire [5:0] lut_237_select = {
                             in_data[4],
                             in_data[37],
                             in_data[16],
                             in_data[40],
                             in_data[3],
                             in_data[24]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [63:0] lut_238_table = 64'b1111000000000000100000000001000011111010000000001111101111110011;
    wire [5:0] lut_238_select = {
                             in_data[60],
                             in_data[17],
                             in_data[56],
                             in_data[15],
                             in_data[55],
                             in_data[45]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [63:0] lut_239_table = 64'b0000001100100011001000110010101100111011001110110011101100111011;
    wire [5:0] lut_239_select = {
                             in_data[46],
                             in_data[29],
                             in_data[58],
                             in_data[38],
                             in_data[26],
                             in_data[11]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [63:0] lut_240_table = 64'b1100110011111111110011001100110011111111111111111100110011000100;
    wire [5:0] lut_240_select = {
                             in_data[28],
                             in_data[22],
                             in_data[20],
                             in_data[61],
                             in_data[51],
                             in_data[23]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [63:0] lut_241_table = 64'b0101000100000000011101110101000101110111000100000111011101010111;
    wire [5:0] lut_241_select = {
                             in_data[25],
                             in_data[47],
                             in_data[29],
                             in_data[58],
                             in_data[63],
                             in_data[4]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [63:0] lut_242_table = 64'b0000111100001100010111110000010100000111000000000011111100000001;
    wire [5:0] lut_242_select = {
                             in_data[1],
                             in_data[0],
                             in_data[35],
                             in_data[41],
                             in_data[18],
                             in_data[7]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [63:0] lut_243_table = 64'b0111011101010011000001000000000011111111111111110100110111111111;
    wire [5:0] lut_243_select = {
                             in_data[56],
                             in_data[52],
                             in_data[13],
                             in_data[32],
                             in_data[2],
                             in_data[39]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [63:0] lut_244_table = 64'b1111011101110111111101110101000111110010001100100111001000110000;
    wire [5:0] lut_244_select = {
                             in_data[44],
                             in_data[10],
                             in_data[57],
                             in_data[33],
                             in_data[42],
                             in_data[15]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [63:0] lut_245_table = 64'b1110101011111010001000001111101010000000101010000000010011101110;
    wire [5:0] lut_245_select = {
                             in_data[31],
                             in_data[50],
                             in_data[59],
                             in_data[55],
                             in_data[5],
                             in_data[38]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [63:0] lut_246_table = 64'b1110111010001000111111101000100011000000100000001111000010000000;
    wire [5:0] lut_246_select = {
                             in_data[14],
                             in_data[8],
                             in_data[26],
                             in_data[12],
                             in_data[53],
                             in_data[19]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [63:0] lut_247_table = 64'b1001111111011111000000001000100010011111100111110000000000001000;
    wire [5:0] lut_247_select = {
                             in_data[40],
                             in_data[16],
                             in_data[48],
                             in_data[60],
                             in_data[27],
                             in_data[17]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [63:0] lut_248_table = 64'b1011001011111111001000001011001010110010111110110010000010110000;
    wire [5:0] lut_248_select = {
                             in_data[46],
                             in_data[24],
                             in_data[11],
                             in_data[45],
                             in_data[62],
                             in_data[6]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [63:0] lut_249_table = 64'b0000000000100010000011111011111100000000001000110000101000111011;
    wire [5:0] lut_249_select = {
                             in_data[21],
                             in_data[30],
                             in_data[43],
                             in_data[3],
                             in_data[36],
                             in_data[37]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [63:0] lut_250_table = 64'b0101010100000000111111110000000011111111010111101111111110001000;
    wire [5:0] lut_250_select = {
                             in_data[61],
                             in_data[4],
                             in_data[54],
                             in_data[49],
                             in_data[34],
                             in_data[9]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [63:0] lut_251_table = 64'b0000000011010101100000001111111100000010111111111000000011111010;
    wire [5:0] lut_251_select = {
                             in_data[10],
                             in_data[15],
                             in_data[8],
                             in_data[50],
                             in_data[37],
                             in_data[16]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [63:0] lut_252_table = 64'b1111111111111110111111111000000011111101111010001111111110000000;
    wire [5:0] lut_252_select = {
                             in_data[33],
                             in_data[28],
                             in_data[29],
                             in_data[12],
                             in_data[41],
                             in_data[26]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [63:0] lut_253_table = 64'b1111101110110011001100110011001011111111111110111111111100010011;
    wire [5:0] lut_253_select = {
                             in_data[30],
                             in_data[58],
                             in_data[48],
                             in_data[23],
                             in_data[11],
                             in_data[13]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [63:0] lut_254_table = 64'b1100000011100000010000000100000011111110111111111111010011110000;
    wire [5:0] lut_254_select = {
                             in_data[59],
                             in_data[35],
                             in_data[39],
                             in_data[3],
                             in_data[63],
                             in_data[55]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [63:0] lut_255_table = 64'b0000010000000100000000000000010001000111110111110000010101010101;
    wire [5:0] lut_255_select = {
                             in_data[47],
                             in_data[0],
                             in_data[24],
                             in_data[18],
                             in_data[57],
                             in_data[43]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [63:0] lut_256_table = 64'b1010101110101010101010101010101010101010100010101010101010101010;
    wire [5:0] lut_256_select = {
                             in_data[27],
                             in_data[7],
                             in_data[21],
                             in_data[62],
                             in_data[38],
                             in_data[32]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [63:0] lut_257_table = 64'b0000100011111110110011111111111100001010101010101010111010101010;
    wire [5:0] lut_257_select = {
                             in_data[20],
                             in_data[1],
                             in_data[5],
                             in_data[44],
                             in_data[36],
                             in_data[56]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [63:0] lut_258_table = 64'b0101000000010001010101010011011111010101010101010101010001010100;
    wire [5:0] lut_258_select = {
                             in_data[51],
                             in_data[45],
                             in_data[46],
                             in_data[14],
                             in_data[6],
                             in_data[42]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [63:0] lut_259_table = 64'b1101111101001100010011110100010011001111000001000100111100000100;
    wire [5:0] lut_259_select = {
                             in_data[60],
                             in_data[22],
                             in_data[40],
                             in_data[53],
                             in_data[31],
                             in_data[19]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [63:0] lut_260_table = 64'b0100010111011111010000000101111100000100010111110000000001011111;
    wire [5:0] lut_260_select = {
                             in_data[35],
                             in_data[28],
                             in_data[52],
                             in_data[25],
                             in_data[17],
                             in_data[2]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [63:0] lut_261_table = 64'b0000000100010111000000010000011100010101000101110001001100110111;
    wire [5:0] lut_261_select = {
                             in_data[14],
                             in_data[46],
                             in_data[12],
                             in_data[27],
                             in_data[33],
                             in_data[55]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [63:0] lut_262_table = 64'b1111111111111011001100100000000011111111111110101010100000000000;
    wire [5:0] lut_262_select = {
                             in_data[49],
                             in_data[10],
                             in_data[38],
                             in_data[3],
                             in_data[30],
                             in_data[18]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [63:0] lut_263_table = 64'b0101110101010010010111110101111100001000000000000000000000001010;
    wire [5:0] lut_263_select = {
                             in_data[63],
                             in_data[31],
                             in_data[16],
                             in_data[54],
                             in_data[37],
                             in_data[45]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [63:0] lut_264_table = 64'b0000010001111101000000010000000000000111111111110011111110111111;
    wire [5:0] lut_264_select = {
                             in_data[32],
                             in_data[40],
                             in_data[43],
                             in_data[60],
                             in_data[48],
                             in_data[61]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [63:0] lut_265_table = 64'b1110010011000100111101100100010011100000000000001111011101000000;
    wire [5:0] lut_265_select = {
                             in_data[5],
                             in_data[57],
                             in_data[26],
                             in_data[44],
                             in_data[41],
                             in_data[11]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [63:0] lut_266_table = 64'b0001000100000000110101011100010001110011001100011111011111110101;
    wire [5:0] lut_266_select = {
                             in_data[6],
                             in_data[15],
                             in_data[21],
                             in_data[39],
                             in_data[1],
                             in_data[51]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [63:0] lut_267_table = 64'b1011110001110000111010001000000010111000111100001010100000000000;
    wire [5:0] lut_267_select = {
                             in_data[29],
                             in_data[13],
                             in_data[53],
                             in_data[7],
                             in_data[62],
                             in_data[19]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [63:0] lut_268_table = 64'b0010101100110011111011110111011100010000000000000101010100000000;
    wire [5:0] lut_268_select = {
                             in_data[36],
                             in_data[47],
                             in_data[50],
                             in_data[4],
                             in_data[8],
                             in_data[56]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [63:0] lut_269_table = 64'b0111011100110111000000000011001100000100001101110000000000100011;
    wire [5:0] lut_269_select = {
                             in_data[59],
                             in_data[34],
                             in_data[42],
                             in_data[24],
                             in_data[0],
                             in_data[22]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [63:0] lut_270_table = 64'b0010001000000000101000101110101010101010101010101010101011111010;
    wire [5:0] lut_270_select = {
                             in_data[14],
                             in_data[32],
                             in_data[20],
                             in_data[23],
                             in_data[58],
                             in_data[9]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [63:0] lut_271_table = 64'b1111111110111111000000010000001101111111111111110101000101010111;
    wire [5:0] lut_271_select = {
                             in_data[41],
                             in_data[25],
                             in_data[46],
                             in_data[48],
                             in_data[47],
                             in_data[42]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [63:0] lut_272_table = 64'b1111111011111111100000001010101010101010111011101010100010101010;
    wire [5:0] lut_272_select = {
                             in_data[18],
                             in_data[38],
                             in_data[60],
                             in_data[15],
                             in_data[12],
                             in_data[43]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [63:0] lut_273_table = 64'b1010001010101000101110101111101100101011001000101011001110111011;
    wire [5:0] lut_273_select = {
                             in_data[11],
                             in_data[29],
                             in_data[37],
                             in_data[4],
                             in_data[55],
                             in_data[19]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [63:0] lut_274_table = 64'b0101000011010000010100000100000011111011111111110101010101010101;
    wire [5:0] lut_274_select = {
                             in_data[45],
                             in_data[21],
                             in_data[49],
                             in_data[36],
                             in_data[54],
                             in_data[33]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [63:0] lut_275_table = 64'b0011001000100010111110111111101000110010111100101111001110111010;
    wire [5:0] lut_275_select = {
                             in_data[40],
                             in_data[3],
                             in_data[17],
                             in_data[22],
                             in_data[26],
                             in_data[27]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [63:0] lut_276_table = 64'b1111001101110011011100110111001101110000000100000000000000010011;
    wire [5:0] lut_276_select = {
                             in_data[7],
                             in_data[61],
                             in_data[16],
                             in_data[57],
                             in_data[31],
                             in_data[53]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [63:0] lut_277_table = 64'b1111001110111011111110111011101101110000000000001111000100110000;
    wire [5:0] lut_277_select = {
                             in_data[6],
                             in_data[28],
                             in_data[39],
                             in_data[30],
                             in_data[10],
                             in_data[8]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [63:0] lut_278_table = 64'b1111111011111110011100110111001000000000000100000001000000000000;
    wire [5:0] lut_278_select = {
                             in_data[5],
                             in_data[34],
                             in_data[59],
                             in_data[51],
                             in_data[35],
                             in_data[56]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [63:0] lut_279_table = 64'b0011000000000000001100000000000011111011001100101111001100110000;
    wire [5:0] lut_279_select = {
                             in_data[44],
                             in_data[62],
                             in_data[50],
                             in_data[2],
                             in_data[24],
                             in_data[1]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [63:0] lut_280_table = 64'b0100111101001111010001010100010101001111010011110000000001000100;
    wire [5:0] lut_280_select = {
                             in_data[8],
                             in_data[30],
                             in_data[63],
                             in_data[52],
                             in_data[0],
                             in_data[13]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [63:0] lut_281_table = 64'b1111111101010101111111110101010101011111010001011101111101010101;
    wire [5:0] lut_281_select = {
                             in_data[42],
                             in_data[43],
                             in_data[19],
                             in_data[53],
                             in_data[7],
                             in_data[22]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [63:0] lut_282_table = 64'b1000101101000110100010110000111110001111110011110000101001001110;
    wire [5:0] lut_282_select = {
                             in_data[20],
                             in_data[2],
                             in_data[5],
                             in_data[3],
                             in_data[16],
                             in_data[1]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [63:0] lut_283_table = 64'b1110000011101100101000001111111000100000111011001010000011111111;
    wire [5:0] lut_283_select = {
                             in_data[49],
                             in_data[41],
                             in_data[24],
                             in_data[14],
                             in_data[59],
                             in_data[29]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [63:0] lut_284_table = 64'b0000101110101011101111111011111100001010101110111011101110111011;
    wire [5:0] lut_284_select = {
                             in_data[39],
                             in_data[37],
                             in_data[18],
                             in_data[12],
                             in_data[48],
                             in_data[31]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [63:0] lut_285_table = 64'b0000101000000000000011100010000000001111000000000110111100001010;
    wire [5:0] lut_285_select = {
                             in_data[62],
                             in_data[56],
                             in_data[9],
                             in_data[38],
                             in_data[10],
                             in_data[47]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [63:0] lut_286_table = 64'b0000000000000000010101010000000011111111111101001111111111110111;
    wire [5:0] lut_286_select = {
                             in_data[44],
                             in_data[36],
                             in_data[15],
                             in_data[4],
                             in_data[46],
                             in_data[25]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [63:0] lut_287_table = 64'b0101000001010000010100001111000011110010111100101111000011111011;
    wire [5:0] lut_287_select = {
                             in_data[60],
                             in_data[33],
                             in_data[58],
                             in_data[61],
                             in_data[40],
                             in_data[26]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [63:0] lut_288_table = 64'b0101111100010101010111110101111101011111000111110001000100010101;
    wire [5:0] lut_288_select = {
                             in_data[23],
                             in_data[51],
                             in_data[17],
                             in_data[6],
                             in_data[11],
                             in_data[32]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [63:0] lut_289_table = 64'b0000000000010101110100011111111100010101000001111111110111111111;
    wire [5:0] lut_289_select = {
                             in_data[34],
                             in_data[54],
                             in_data[55],
                             in_data[27],
                             in_data[50],
                             in_data[57]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [63:0] lut_290_table = 64'b0000000000001010000000000010111100101010101111111011101111111111;
    wire [5:0] lut_290_select = {
                             in_data[14],
                             in_data[44],
                             in_data[28],
                             in_data[35],
                             in_data[45],
                             in_data[21]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [63:0] lut_291_table = 64'b1100010011111111010011101111111100000000011100110010000011110111;
    wire [5:0] lut_291_select = {
                             in_data[25],
                             in_data[58],
                             in_data[52],
                             in_data[63],
                             in_data[3],
                             in_data[19]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [63:0] lut_292_table = 64'b1111111100011111101111110000111000110011000001011011111100001111;
    wire [5:0] lut_292_select = {
                             in_data[57],
                             in_data[38],
                             in_data[36],
                             in_data[17],
                             in_data[33],
                             in_data[4]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [63:0] lut_293_table = 64'b0000010000000000110111110000000001000100000000001111111111111101;
    wire [5:0] lut_293_select = {
                             in_data[29],
                             in_data[24],
                             in_data[32],
                             in_data[42],
                             in_data[11],
                             in_data[59]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [63:0] lut_294_table = 64'b1110110000000000111111000000000011111111100010001111111100001100;
    wire [5:0] lut_294_select = {
                             in_data[6],
                             in_data[31],
                             in_data[2],
                             in_data[23],
                             in_data[55],
                             in_data[47]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [63:0] lut_295_table = 64'b1100110000001101110111010100111111011111000011111111111101011111;
    wire [5:0] lut_295_select = {
                             in_data[18],
                             in_data[50],
                             in_data[53],
                             in_data[27],
                             in_data[16],
                             in_data[40]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [63:0] lut_296_table = 64'b0011001100000000101110110000000011110011101100001111001100000000;
    wire [5:0] lut_296_select = {
                             in_data[39],
                             in_data[49],
                             in_data[37],
                             in_data[0],
                             in_data[41],
                             in_data[10]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [63:0] lut_297_table = 64'b1010110010101000100010001000100011001111111011111100111010101110;
    wire [5:0] lut_297_select = {
                             in_data[15],
                             in_data[61],
                             in_data[12],
                             in_data[5],
                             in_data[56],
                             in_data[62]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [63:0] lut_298_table = 64'b0000010100001111000001010000000000001111000011110000111100001111;
    wire [5:0] lut_298_select = {
                             in_data[22],
                             in_data[20],
                             in_data[7],
                             in_data[51],
                             in_data[30],
                             in_data[9]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [63:0] lut_299_table = 64'b1111010011110101011000001111010111000000111101000111000011110001;
    wire [5:0] lut_299_select = {
                             in_data[43],
                             in_data[48],
                             in_data[34],
                             in_data[1],
                             in_data[60],
                             in_data[13]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [63:0] lut_300_table = 64'b1110111111001111111011111100111011001111000001001000111000001100;
    wire [5:0] lut_300_select = {
                             in_data[42],
                             in_data[21],
                             in_data[54],
                             in_data[8],
                             in_data[26],
                             in_data[46]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [63:0] lut_301_table = 64'b0111111111111111001100110011101111101111111111110010111100101110;
    wire [5:0] lut_301_select = {
                             in_data[10],
                             in_data[25],
                             in_data[57],
                             in_data[48],
                             in_data[56],
                             in_data[53]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [63:0] lut_302_table = 64'b0100010001001100010001000100010001000100010011100100000001011110;
    wire [5:0] lut_302_select = {
                             in_data[36],
                             in_data[7],
                             in_data[11],
                             in_data[63],
                             in_data[30],
                             in_data[4]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [63:0] lut_303_table = 64'b0000100011101110000000001000111010001111111011110011111110101111;
    wire [5:0] lut_303_select = {
                             in_data[1],
                             in_data[17],
                             in_data[61],
                             in_data[58],
                             in_data[33],
                             in_data[24]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [63:0] lut_304_table = 64'b1010101010101010101110100010101010101010101010101011001000111011;
    wire [5:0] lut_304_select = {
                             in_data[50],
                             in_data[27],
                             in_data[28],
                             in_data[62],
                             in_data[35],
                             in_data[22]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [63:0] lut_305_table = 64'b0000100010101010000010001010101000001110101011111010111010101110;
    wire [5:0] lut_305_select = {
                             in_data[31],
                             in_data[47],
                             in_data[41],
                             in_data[38],
                             in_data[12],
                             in_data[13]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [63:0] lut_306_table = 64'b0000010001011101010011000101111101000000010101010101010011011101;
    wire [5:0] lut_306_select = {
                             in_data[16],
                             in_data[49],
                             in_data[5],
                             in_data[32],
                             in_data[2],
                             in_data[44]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [63:0] lut_307_table = 64'b1111000101110001111111110111011101110000010100001111011101010001;
    wire [5:0] lut_307_select = {
                             in_data[51],
                             in_data[45],
                             in_data[0],
                             in_data[52],
                             in_data[39],
                             in_data[37]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [63:0] lut_308_table = 64'b1100111100000000100001000000000011101111000000001100110010000000;
    wire [5:0] lut_308_select = {
                             in_data[60],
                             in_data[43],
                             in_data[19],
                             in_data[40],
                             in_data[3],
                             in_data[23]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [63:0] lut_309_table = 64'b0000111110001111010001111101111111001111100011110000110100001101;
    wire [5:0] lut_309_select = {
                             in_data[20],
                             in_data[9],
                             in_data[14],
                             in_data[6],
                             in_data[15],
                             in_data[29]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [63:0] lut_310_table = 64'b0011001100110001001110111111010100110011001100001011101101110000;
    wire [5:0] lut_310_select = {
                             in_data[54],
                             in_data[62],
                             in_data[34],
                             in_data[55],
                             in_data[18],
                             in_data[59]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [63:0] lut_311_table = 64'b1110111110001010101011101000100011101110101010001110101010101000;
    wire [5:0] lut_311_select = {
                             in_data[27],
                             in_data[47],
                             in_data[28],
                             in_data[22],
                             in_data[38],
                             in_data[14]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [63:0] lut_312_table = 64'b0101000001110001011100011111011101010000110100010101010101110111;
    wire [5:0] lut_312_select = {
                             in_data[46],
                             in_data[3],
                             in_data[23],
                             in_data[12],
                             in_data[17],
                             in_data[33]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [63:0] lut_313_table = 64'b1101010100010101010101010101010111110101010101011101010101010101;
    wire [5:0] lut_313_select = {
                             in_data[20],
                             in_data[58],
                             in_data[40],
                             in_data[42],
                             in_data[26],
                             in_data[41]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [63:0] lut_314_table = 64'b0010101000100010001011100011101000111111001100100000101100100010;
    wire [5:0] lut_314_select = {
                             in_data[53],
                             in_data[1],
                             in_data[0],
                             in_data[60],
                             in_data[5],
                             in_data[21]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [63:0] lut_315_table = 64'b0000000100000000000100010000000000011101111111110001011100111111;
    wire [5:0] lut_315_select = {
                             in_data[4],
                             in_data[48],
                             in_data[11],
                             in_data[16],
                             in_data[43],
                             in_data[24]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [63:0] lut_316_table = 64'b0001000110110000000100000101000011110001111100110101000011110001;
    wire [5:0] lut_316_select = {
                             in_data[57],
                             in_data[63],
                             in_data[6],
                             in_data[50],
                             in_data[36],
                             in_data[31]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [63:0] lut_317_table = 64'b1111111110110011001111110011111111100000101000001011111110101111;
    wire [5:0] lut_317_select = {
                             in_data[51],
                             in_data[56],
                             in_data[25],
                             in_data[7],
                             in_data[10],
                             in_data[9]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [63:0] lut_318_table = 64'b0000000001000100010101111111110100000000010001000001111111010110;
    wire [5:0] lut_318_select = {
                             in_data[44],
                             in_data[45],
                             in_data[35],
                             in_data[19],
                             in_data[8],
                             in_data[30]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [63:0] lut_319_table = 64'b1010101010101010101010101110101000101010001010101010101110101010;
    wire [5:0] lut_319_select = {
                             in_data[13],
                             in_data[32],
                             in_data[29],
                             in_data[61],
                             in_data[39],
                             in_data[2]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [63:0] lut_320_table = 64'b0011111100000000001111110000101010101111000000001011111100000010;
    wire [5:0] lut_320_select = {
                             in_data[39],
                             in_data[57],
                             in_data[49],
                             in_data[37],
                             in_data[52],
                             in_data[15]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [63:0] lut_321_table = 64'b0011011100110111000101110001001100010011001111110111011101111111;
    wire [5:0] lut_321_select = {
                             in_data[26],
                             in_data[8],
                             in_data[1],
                             in_data[17],
                             in_data[20],
                             in_data[12]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [63:0] lut_322_table = 64'b0000000011111000101010101111111000000000111100000000001011111000;
    wire [5:0] lut_322_select = {
                             in_data[16],
                             in_data[22],
                             in_data[50],
                             in_data[53],
                             in_data[63],
                             in_data[43]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [63:0] lut_323_table = 64'b1111000011111110001000001111111011111000111111101100000011111110;
    wire [5:0] lut_323_select = {
                             in_data[46],
                             in_data[4],
                             in_data[48],
                             in_data[31],
                             in_data[3],
                             in_data[47]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [63:0] lut_324_table = 64'b0000000111111010110111111111111100000001000110110101111111111101;
    wire [5:0] lut_324_select = {
                             in_data[19],
                             in_data[36],
                             in_data[28],
                             in_data[29],
                             in_data[34],
                             in_data[62]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [63:0] lut_325_table = 64'b0000001000001000100000000000100010101010111011101110111011101110;
    wire [5:0] lut_325_select = {
                             in_data[18],
                             in_data[6],
                             in_data[61],
                             in_data[0],
                             in_data[56],
                             in_data[42]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [63:0] lut_326_table = 64'b1111100111111001111110111111111100000000000000000010001100100010;
    wire [5:0] lut_326_select = {
                             in_data[38],
                             in_data[44],
                             in_data[45],
                             in_data[10],
                             in_data[25],
                             in_data[13]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [63:0] lut_327_table = 64'b0000010100000111000010100000001111101111111011111111111111101111;
    wire [5:0] lut_327_select = {
                             in_data[27],
                             in_data[54],
                             in_data[32],
                             in_data[59],
                             in_data[5],
                             in_data[14]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [63:0] lut_328_table = 64'b0000101010101010110010101110111000000000000000001100100001000000;
    wire [5:0] lut_328_select = {
                             in_data[33],
                             in_data[55],
                             in_data[23],
                             in_data[41],
                             in_data[9],
                             in_data[11]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [63:0] lut_329_table = 64'b0011001100110111000000100011001101110011011111110011001101110011;
    wire [5:0] lut_329_select = {
                             in_data[7],
                             in_data[30],
                             in_data[58],
                             in_data[51],
                             in_data[2],
                             in_data[60]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [63:0] lut_330_table = 64'b1111111111111111001101110001010100110000000100010011001100110011;
    wire [5:0] lut_330_select = {
                             in_data[12],
                             in_data[19],
                             in_data[24],
                             in_data[40],
                             in_data[21],
                             in_data[35]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [63:0] lut_331_table = 64'b1001111100011011000010110000101111111111101111111001111100101011;
    wire [5:0] lut_331_select = {
                             in_data[63],
                             in_data[56],
                             in_data[58],
                             in_data[22],
                             in_data[25],
                             in_data[48]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [63:0] lut_332_table = 64'b0010101010101010111111111111111100000000000000001111101011001100;
    wire [5:0] lut_332_select = {
                             in_data[54],
                             in_data[26],
                             in_data[42],
                             in_data[4],
                             in_data[44],
                             in_data[51]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [63:0] lut_333_table = 64'b1011000111111111001000001111010010111011111111110010001111110111;
    wire [5:0] lut_333_select = {
                             in_data[32],
                             in_data[39],
                             in_data[47],
                             in_data[34],
                             in_data[45],
                             in_data[41]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [63:0] lut_334_table = 64'b0000000001011101000101000101110100000100010111010101010101011111;
    wire [5:0] lut_334_select = {
                             in_data[30],
                             in_data[23],
                             in_data[29],
                             in_data[38],
                             in_data[8],
                             in_data[60]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [63:0] lut_335_table = 64'b1010000000100000111101001111110100100000001000001010000000100100;
    wire [5:0] lut_335_select = {
                             in_data[17],
                             in_data[36],
                             in_data[62],
                             in_data[20],
                             in_data[15],
                             in_data[43]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [63:0] lut_336_table = 64'b0000000100000001000000000000100000001101000011011100111111111111;
    wire [5:0] lut_336_select = {
                             in_data[57],
                             in_data[59],
                             in_data[16],
                             in_data[13],
                             in_data[3],
                             in_data[49]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [63:0] lut_337_table = 64'b1011001100110010001100110010000000110011001100110011001100110001;
    wire [5:0] lut_337_select = {
                             in_data[50],
                             in_data[37],
                             in_data[1],
                             in_data[33],
                             in_data[28],
                             in_data[52]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [63:0] lut_338_table = 64'b1010001011111111001100101111111100000000001100110000000001110111;
    wire [5:0] lut_338_select = {
                             in_data[14],
                             in_data[31],
                             in_data[27],
                             in_data[18],
                             in_data[0],
                             in_data[5]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [63:0] lut_339_table = 64'b1110000011100000111110101111101011010000110100001111000011110010;
    wire [5:0] lut_339_select = {
                             in_data[53],
                             in_data[55],
                             in_data[10],
                             in_data[6],
                             in_data[61],
                             in_data[2]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [63:0] lut_340_table = 64'b0000101000000011010110110000001000011011000000100101111000001010;
    wire [5:0] lut_340_select = {
                             in_data[4],
                             in_data[8],
                             in_data[46],
                             in_data[7],
                             in_data[11],
                             in_data[9]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [63:0] lut_341_table = 64'b0001000000011101000100000001000000111011111111110111001101111111;
    wire [5:0] lut_341_select = {
                             in_data[36],
                             in_data[58],
                             in_data[55],
                             in_data[12],
                             in_data[38],
                             in_data[22]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [63:0] lut_342_table = 64'b0101110111111111000001010101010100000101010101010000000000000000;
    wire [5:0] lut_342_select = {
                             in_data[42],
                             in_data[21],
                             in_data[20],
                             in_data[60],
                             in_data[52],
                             in_data[33]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [63:0] lut_343_table = 64'b1111001100110010101100100010001000110001000000000000000000000000;
    wire [5:0] lut_343_select = {
                             in_data[1],
                             in_data[48],
                             in_data[56],
                             in_data[41],
                             in_data[16],
                             in_data[0]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [63:0] lut_344_table = 64'b0000100010101111101010101011111100000000000010100000001010111011;
    wire [5:0] lut_344_select = {
                             in_data[34],
                             in_data[39],
                             in_data[5],
                             in_data[63],
                             in_data[14],
                             in_data[50]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [63:0] lut_345_table = 64'b1111110111011101110101011111110101000101010001000101000001010101;
    wire [5:0] lut_345_select = {
                             in_data[23],
                             in_data[53],
                             in_data[57],
                             in_data[43],
                             in_data[10],
                             in_data[30]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [63:0] lut_346_table = 64'b1111110101011101111100001111010010111101010000001111000001000000;
    wire [5:0] lut_346_select = {
                             in_data[47],
                             in_data[32],
                             in_data[15],
                             in_data[29],
                             in_data[18],
                             in_data[25]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [63:0] lut_347_table = 64'b0000110111001100000011001000110000011101111111010000110100001100;
    wire [5:0] lut_347_select = {
                             in_data[26],
                             in_data[44],
                             in_data[28],
                             in_data[62],
                             in_data[45],
                             in_data[3]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [63:0] lut_348_table = 64'b0010001010111011011100111111101110111011101110111111101100110011;
    wire [5:0] lut_348_select = {
                             in_data[6],
                             in_data[31],
                             in_data[17],
                             in_data[27],
                             in_data[24],
                             in_data[49]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [63:0] lut_349_table = 64'b1111110101010000111101010101000011110101011101001111010101010100;
    wire [5:0] lut_349_select = {
                             in_data[40],
                             in_data[59],
                             in_data[37],
                             in_data[51],
                             in_data[61],
                             in_data[19]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [63:0] lut_350_table = 64'b1110101000000010111010001111111010000010000000011111111011111111;
    wire [5:0] lut_350_select = {
                             in_data[49],
                             in_data[37],
                             in_data[2],
                             in_data[54],
                             in_data[13],
                             in_data[35]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [63:0] lut_351_table = 64'b1011001001000000001100110101010101010000010100000101000101010101;
    wire [5:0] lut_351_select = {
                             in_data[22],
                             in_data[38],
                             in_data[27],
                             in_data[10],
                             in_data[46],
                             in_data[63]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [63:0] lut_352_table = 64'b1111110011111000111111111010000011110000111000001111110010000000;
    wire [5:0] lut_352_select = {
                             in_data[55],
                             in_data[58],
                             in_data[41],
                             in_data[14],
                             in_data[24],
                             in_data[48]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [63:0] lut_353_table = 64'b1111111111111111011101110101011101110011010101010011000100010101;
    wire [5:0] lut_353_select = {
                             in_data[8],
                             in_data[20],
                             in_data[6],
                             in_data[36],
                             in_data[17],
                             in_data[33]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [63:0] lut_354_table = 64'b1110111100001111111111111111111100000000000000001111111110011111;
    wire [5:0] lut_354_select = {
                             in_data[51],
                             in_data[19],
                             in_data[32],
                             in_data[15],
                             in_data[28],
                             in_data[50]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [63:0] lut_355_table = 64'b1111110111010100110111000100010011010100010001000100010001000000;
    wire [5:0] lut_355_select = {
                             in_data[21],
                             in_data[43],
                             in_data[39],
                             in_data[53],
                             in_data[7],
                             in_data[9]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [63:0] lut_356_table = 64'b1101111110001100000010100000101011111111100011100000111100000000;
    wire [5:0] lut_356_select = {
                             in_data[52],
                             in_data[59],
                             in_data[23],
                             in_data[30],
                             in_data[56],
                             in_data[18]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [63:0] lut_357_table = 64'b1100010011011101110011001101110101000000110011001100110011011101;
    wire [5:0] lut_357_select = {
                             in_data[26],
                             in_data[34],
                             in_data[1],
                             in_data[61],
                             in_data[12],
                             in_data[44]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [63:0] lut_358_table = 64'b1111101111111011111100001110001010101000101010101010000010101000;
    wire [5:0] lut_358_select = {
                             in_data[45],
                             in_data[11],
                             in_data[40],
                             in_data[57],
                             in_data[62],
                             in_data[5]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [63:0] lut_359_table = 64'b1111101000000000111111111111101000000000000000001101110001110010;
    wire [5:0] lut_359_select = {
                             in_data[29],
                             in_data[25],
                             in_data[0],
                             in_data[42],
                             in_data[3],
                             in_data[16]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub4
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        359:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [         59:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub4_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub4_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub4_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [359:0]  in_data,
            output wire [59:0]  out_data
        );
    
    
    // LUT : 0
    wire [63:0] lut_0_table = 64'b1100110000000000111111111111110111000000000000001111110011010100;
    wire [5:0] lut_0_select = {
                             in_data[111],
                             in_data[82],
                             in_data[280],
                             in_data[316],
                             in_data[302],
                             in_data[8]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [63:0] lut_1_table = 64'b1110111110001010100011101000101011101111100010101000101010001000;
    wire [5:0] lut_1_select = {
                             in_data[20],
                             in_data[289],
                             in_data[203],
                             in_data[344],
                             in_data[191],
                             in_data[73]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [63:0] lut_2_table = 64'b1111101011111010101110100010001011111010001100101011101000100010;
    wire [5:0] lut_2_select = {
                             in_data[310],
                             in_data[148],
                             in_data[47],
                             in_data[10],
                             in_data[278],
                             in_data[71]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [63:0] lut_3_table = 64'b1000100000001000101010101000101011000100000011001100011011001111;
    wire [5:0] lut_3_select = {
                             in_data[330],
                             in_data[120],
                             in_data[98],
                             in_data[178],
                             in_data[44],
                             in_data[133]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [63:0] lut_4_table = 64'b1011001100111011001100110010001100110011001100110011001000000000;
    wire [5:0] lut_4_select = {
                             in_data[132],
                             in_data[234],
                             in_data[48],
                             in_data[129],
                             in_data[259],
                             in_data[334]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [63:0] lut_5_table = 64'b1111111101010111111111110001000101011111000100010000000111000001;
    wire [5:0] lut_5_select = {
                             in_data[0],
                             in_data[65],
                             in_data[30],
                             in_data[193],
                             in_data[298],
                             in_data[41]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [63:0] lut_6_table = 64'b1101000011010100000000000000000011110101111101110111010111111111;
    wire [5:0] lut_6_select = {
                             in_data[206],
                             in_data[359],
                             in_data[347],
                             in_data[40],
                             in_data[135],
                             in_data[205]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [63:0] lut_7_table = 64'b0100010000001101110111011000110100000100110101001101110111111101;
    wire [5:0] lut_7_select = {
                             in_data[338],
                             in_data[341],
                             in_data[61],
                             in_data[254],
                             in_data[320],
                             in_data[275]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [63:0] lut_8_table = 64'b1111010111010100110100011100000011010001111101001101000111010000;
    wire [5:0] lut_8_select = {
                             in_data[200],
                             in_data[101],
                             in_data[194],
                             in_data[274],
                             in_data[78],
                             in_data[329]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [63:0] lut_9_table = 64'b0001011101111111000101111111111100000011000101110000001100111111;
    wire [5:0] lut_9_select = {
                             in_data[157],
                             in_data[322],
                             in_data[265],
                             in_data[327],
                             in_data[141],
                             in_data[355]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [63:0] lut_10_table = 64'b1111111101110000111101110111000001110011001100100011001000100010;
    wire [5:0] lut_10_select = {
                             in_data[218],
                             in_data[235],
                             in_data[252],
                             in_data[37],
                             in_data[36],
                             in_data[296]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [63:0] lut_11_table = 64'b1101010011011101010000001100010011111100111111111101010011111101;
    wire [5:0] lut_11_select = {
                             in_data[125],
                             in_data[159],
                             in_data[124],
                             in_data[32],
                             in_data[53],
                             in_data[224]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [63:0] lut_12_table = 64'b0101111101011111001100111111111100000011000101110000000100010111;
    wire [5:0] lut_12_select = {
                             in_data[123],
                             in_data[147],
                             in_data[340],
                             in_data[115],
                             in_data[171],
                             in_data[96]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [63:0] lut_13_table = 64'b1011001110110010111110111111101110110010001000001111101111110010;
    wire [5:0] lut_13_select = {
                             in_data[181],
                             in_data[222],
                             in_data[263],
                             in_data[168],
                             in_data[128],
                             in_data[232]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [63:0] lut_14_table = 64'b0000010000000000110011010010010000001101000001001101111101001101;
    wire [5:0] lut_14_select = {
                             in_data[293],
                             in_data[276],
                             in_data[352],
                             in_data[104],
                             in_data[19],
                             in_data[94]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [63:0] lut_15_table = 64'b1111000101110001111111110111011101010001000000001111011101010001;
    wire [5:0] lut_15_select = {
                             in_data[144],
                             in_data[79],
                             in_data[267],
                             in_data[272],
                             in_data[317],
                             in_data[112]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [63:0] lut_16_table = 64'b0000010001010101111001010111111100000000000001010000110101011111;
    wire [5:0] lut_16_select = {
                             in_data[353],
                             in_data[116],
                             in_data[337],
                             in_data[58],
                             in_data[97],
                             in_data[247]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [63:0] lut_17_table = 64'b0000111111001111000011100000111010001010110011100000100011001000;
    wire [5:0] lut_17_select = {
                             in_data[304],
                             in_data[221],
                             in_data[182],
                             in_data[34],
                             in_data[319],
                             in_data[77]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [63:0] lut_18_table = 64'b0001001100110011000000010001001100110011101110110001001100111111;
    wire [5:0] lut_18_select = {
                             in_data[152],
                             in_data[216],
                             in_data[33],
                             in_data[167],
                             in_data[291],
                             in_data[339]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [63:0] lut_19_table = 64'b0010111100111011000010110011111100001011101111110000000000001011;
    wire [5:0] lut_19_select = {
                             in_data[74],
                             in_data[45],
                             in_data[315],
                             in_data[4],
                             in_data[220],
                             in_data[166]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [63:0] lut_20_table = 64'b1010000011110010101000001110100011111010111111111010001011111010;
    wire [5:0] lut_20_select = {
                             in_data[64],
                             in_data[266],
                             in_data[262],
                             in_data[312],
                             in_data[172],
                             in_data[21]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [63:0] lut_21_table = 64'b0001000011110011001100000011001111111011111111111010101000111011;
    wire [5:0] lut_21_select = {
                             in_data[54],
                             in_data[311],
                             in_data[211],
                             in_data[51],
                             in_data[26],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [63:0] lut_22_table = 64'b0101000000010000011101010111000011111101001100101111111111110111;
    wire [5:0] lut_22_select = {
                             in_data[43],
                             in_data[107],
                             in_data[1],
                             in_data[52],
                             in_data[332],
                             in_data[118]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [63:0] lut_23_table = 64'b0000001100101011000000000000001000101011101111110000000010101011;
    wire [5:0] lut_23_select = {
                             in_data[202],
                             in_data[188],
                             in_data[195],
                             in_data[335],
                             in_data[49],
                             in_data[35]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [63:0] lut_24_table = 64'b1000000011111000110101001111110111110100111111001101010011111101;
    wire [5:0] lut_24_select = {
                             in_data[17],
                             in_data[155],
                             in_data[270],
                             in_data[241],
                             in_data[149],
                             in_data[269]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [63:0] lut_25_table = 64'b0000111100111111000010000000101011111111111111111000111010101111;
    wire [5:0] lut_25_select = {
                             in_data[63],
                             in_data[69],
                             in_data[248],
                             in_data[142],
                             in_data[176],
                             in_data[357]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [63:0] lut_26_table = 64'b1111111110110010101100100010000011110010001000000010000000000000;
    wire [5:0] lut_26_select = {
                             in_data[231],
                             in_data[236],
                             in_data[324],
                             in_data[11],
                             in_data[179],
                             in_data[131]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [63:0] lut_27_table = 64'b1000010000000000010011010100010111000101010101010101111101011111;
    wire [5:0] lut_27_select = {
                             in_data[16],
                             in_data[164],
                             in_data[256],
                             in_data[223],
                             in_data[122],
                             in_data[86]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [63:0] lut_28_table = 64'b0101000011010101010100001111111101000000110100000101000011110101;
    wire [5:0] lut_28_select = {
                             in_data[80],
                             in_data[346],
                             in_data[84],
                             in_data[244],
                             in_data[2],
                             in_data[283]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [63:0] lut_29_table = 64'b0000001010101011000000000101001110111011111111111011111111111111;
    wire [5:0] lut_29_select = {
                             in_data[264],
                             in_data[130],
                             in_data[186],
                             in_data[249],
                             in_data[42],
                             in_data[331]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [63:0] lut_30_table = 64'b0011001101110100001100100011011000000001000101110000000000000001;
    wire [5:0] lut_30_select = {
                             in_data[286],
                             in_data[99],
                             in_data[284],
                             in_data[333],
                             in_data[151],
                             in_data[321]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [63:0] lut_31_table = 64'b0000000000010000010101010111000100100000001100110111010111100010;
    wire [5:0] lut_31_select = {
                             in_data[228],
                             in_data[67],
                             in_data[160],
                             in_data[3],
                             in_data[189],
                             in_data[243]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [63:0] lut_32_table = 64'b0000110100001111000011000000000011111111000111110001111100000011;
    wire [5:0] lut_32_select = {
                             in_data[60],
                             in_data[62],
                             in_data[294],
                             in_data[198],
                             in_data[229],
                             in_data[309]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [63:0] lut_33_table = 64'b0000101000000000001110110010001110101010000000001011100000000000;
    wire [5:0] lut_33_select = {
                             in_data[214],
                             in_data[100],
                             in_data[318],
                             in_data[207],
                             in_data[204],
                             in_data[39]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [63:0] lut_34_table = 64'b1110111011101110000000001110000011111110111011101110100011111010;
    wire [5:0] lut_34_select = {
                             in_data[292],
                             in_data[279],
                             in_data[76],
                             in_data[81],
                             in_data[197],
                             in_data[113]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [63:0] lut_35_table = 64'b0000000001010000010100001111111101010000010100000101000011111101;
    wire [5:0] lut_35_select = {
                             in_data[190],
                             in_data[14],
                             in_data[209],
                             in_data[177],
                             in_data[92],
                             in_data[314]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [63:0] lut_36_table = 64'b0011000101110001011101110111011100010000000100000111000100010001;
    wire [5:0] lut_36_select = {
                             in_data[240],
                             in_data[27],
                             in_data[290],
                             in_data[136],
                             in_data[287],
                             in_data[273]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [63:0] lut_37_table = 64'b0100110011011101000000000100110111011101111111010100110011011100;
    wire [5:0] lut_37_select = {
                             in_data[22],
                             in_data[46],
                             in_data[102],
                             in_data[323],
                             in_data[351],
                             in_data[134]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [63:0] lut_38_table = 64'b1111010101110000010100000101000011111111111100011111000101110000;
    wire [5:0] lut_38_select = {
                             in_data[119],
                             in_data[251],
                             in_data[169],
                             in_data[183],
                             in_data[162],
                             in_data[108]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [63:0] lut_39_table = 64'b0000000100010111000111110111111100000001000111010001111111011111;
    wire [5:0] lut_39_select = {
                             in_data[253],
                             in_data[215],
                             in_data[114],
                             in_data[28],
                             in_data[336],
                             in_data[328]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [63:0] lut_40_table = 64'b1100010011000100111011111100111010001110000010001110111111001110;
    wire [5:0] lut_40_select = {
                             in_data[75],
                             in_data[173],
                             in_data[326],
                             in_data[127],
                             in_data[5],
                             in_data[25]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [63:0] lut_41_table = 64'b0000010101001100010111110100111101000100110011001100110111011111;
    wire [5:0] lut_41_select = {
                             in_data[210],
                             in_data[68],
                             in_data[225],
                             in_data[12],
                             in_data[345],
                             in_data[174]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [63:0] lut_42_table = 64'b1011101000100000101110111011101010110010000000001011101110111010;
    wire [5:0] lut_42_select = {
                             in_data[238],
                             in_data[139],
                             in_data[93],
                             in_data[175],
                             in_data[89],
                             in_data[230]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [63:0] lut_43_table = 64'b1111101111111011101000101011101000110010101100110000000000110011;
    wire [5:0] lut_43_select = {
                             in_data[271],
                             in_data[138],
                             in_data[105],
                             in_data[307],
                             in_data[66],
                             in_data[91]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [63:0] lut_44_table = 64'b0000010000000000010011010000110011001101010011001101111111001111;
    wire [5:0] lut_44_select = {
                             in_data[150],
                             in_data[90],
                             in_data[301],
                             in_data[233],
                             in_data[95],
                             in_data[137]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [63:0] lut_45_table = 64'b0111110100000000010111110000110111011101000000001101111111001101;
    wire [5:0] lut_45_select = {
                             in_data[260],
                             in_data[59],
                             in_data[145],
                             in_data[308],
                             in_data[299],
                             in_data[13]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [63:0] lut_46_table = 64'b1000111011101111100011101110111100000000100011100000100011001111;
    wire [5:0] lut_46_select = {
                             in_data[226],
                             in_data[170],
                             in_data[250],
                             in_data[354],
                             in_data[261],
                             in_data[121]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [63:0] lut_47_table = 64'b1111110100000000001100000000000011111111101100000011000000110000;
    wire [5:0] lut_47_select = {
                             in_data[297],
                             in_data[70],
                             in_data[285],
                             in_data[288],
                             in_data[180],
                             in_data[83]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [63:0] lut_48_table = 64'b0010101000000010001010110010101000101110001110101111111110111011;
    wire [5:0] lut_48_select = {
                             in_data[55],
                             in_data[184],
                             in_data[117],
                             in_data[303],
                             in_data[245],
                             in_data[349]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [63:0] lut_49_table = 64'b1010111110101111001101111010001100011111000000110000000000000000;
    wire [5:0] lut_49_select = {
                             in_data[246],
                             in_data[161],
                             in_data[163],
                             in_data[50],
                             in_data[140],
                             in_data[56]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [63:0] lut_50_table = 64'b0111000101110000111101111110001001010000010000001111010101110000;
    wire [5:0] lut_50_select = {
                             in_data[306],
                             in_data[356],
                             in_data[277],
                             in_data[268],
                             in_data[358],
                             in_data[109]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [63:0] lut_51_table = 64'b1111111100010111010101110000000111111100011101110111111100000001;
    wire [5:0] lut_51_select = {
                             in_data[219],
                             in_data[213],
                             in_data[305],
                             in_data[9],
                             in_data[143],
                             in_data[199]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [63:0] lut_52_table = 64'b1010000010000000101110111010001010111000101000001111101110111010;
    wire [5:0] lut_52_select = {
                             in_data[165],
                             in_data[154],
                             in_data[126],
                             in_data[87],
                             in_data[31],
                             in_data[342]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [63:0] lut_53_table = 64'b1000100010001000111010001010100010001000100010001111111011101100;
    wire [5:0] lut_53_select = {
                             in_data[7],
                             in_data[153],
                             in_data[300],
                             in_data[212],
                             in_data[281],
                             in_data[192]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [63:0] lut_54_table = 64'b0000101000001010110011101100110010001110101011101111111111101111;
    wire [5:0] lut_54_select = {
                             in_data[23],
                             in_data[313],
                             in_data[239],
                             in_data[6],
                             in_data[110],
                             in_data[29]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [63:0] lut_55_table = 64'b0000000000000001000000110001001100000111000101110111011101111111;
    wire [5:0] lut_55_select = {
                             in_data[255],
                             in_data[15],
                             in_data[227],
                             in_data[85],
                             in_data[18],
                             in_data[196]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [63:0] lut_56_table = 64'b0100000011011100010000001100010011111100111111011101010011110000;
    wire [5:0] lut_56_select = {
                             in_data[38],
                             in_data[217],
                             in_data[106],
                             in_data[103],
                             in_data[57],
                             in_data[24]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [63:0] lut_57_table = 64'b0000000001000000010001001101110100000000111101001100010011111101;
    wire [5:0] lut_57_select = {
                             in_data[237],
                             in_data[146],
                             in_data[156],
                             in_data[242],
                             in_data[282],
                             in_data[257]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [63:0] lut_58_table = 64'b1011001011111011001000001010000010101011101110111010100011101010;
    wire [5:0] lut_58_select = {
                             in_data[185],
                             in_data[158],
                             in_data[350],
                             in_data[343],
                             in_data[325],
                             in_data[88]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [63:0] lut_59_table = 64'b0011010100100001011111110111010100000000000000000101010100000101;
    wire [5:0] lut_59_select = {
                             in_data[72],
                             in_data[295],
                             in_data[258],
                             in_data[187],
                             in_data[348],
                             in_data[201]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub5
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [         59:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [          9:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub5_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub5_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub5_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [59:0]  in_data,
            output wire [9:0]  out_data
        );
    
    
    // LUT : 0
    wire [63:0] lut_0_table = 64'b0000000000000000000000000001000000000000000000000000000001010000;
    wire [5:0] lut_0_select = {
                             in_data[33],
                             in_data[52],
                             in_data[32],
                             in_data[27],
                             in_data[17],
                             in_data[8]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [63:0] lut_1_table = 64'b0001000000010000000000000000000001110001010100000000000000000000;
    wire [5:0] lut_1_select = {
                             in_data[20],
                             in_data[53],
                             in_data[14],
                             in_data[26],
                             in_data[25],
                             in_data[51]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [63:0] lut_2_table = 64'b0000000000100000000000000000000010100000101100100000000000100010;
    wire [5:0] lut_2_select = {
                             in_data[57],
                             in_data[16],
                             in_data[47],
                             in_data[10],
                             in_data[3],
                             in_data[24]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [63:0] lut_3_table = 64'b0000000011001000000000001000000011001000111011000000000010001000;
    wire [5:0] lut_3_select = {
                             in_data[37],
                             in_data[21],
                             in_data[58],
                             in_data[22],
                             in_data[44],
                             in_data[19]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [63:0] lut_4_table = 64'b0001000000010000011101010001000100000000000000000001000100010000;
    wire [5:0] lut_4_select = {
                             in_data[45],
                             in_data[31],
                             in_data[48],
                             in_data[9],
                             in_data[7],
                             in_data[15]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [63:0] lut_5_table = 64'b0000000000001000000000000000000000001010100011110000100000001010;
    wire [5:0] lut_5_select = {
                             in_data[0],
                             in_data[28],
                             in_data[30],
                             in_data[34],
                             in_data[2],
                             in_data[41]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [63:0] lut_6_table = 64'b0100010000000000000000000000000001001101000001000000000000000000;
    wire [5:0] lut_6_select = {
                             in_data[18],
                             in_data[54],
                             in_data[35],
                             in_data[40],
                             in_data[1],
                             in_data[50]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [63:0] lut_7_table = 64'b0000000000000000000000000000000001000101000001010000010100000000;
    wire [5:0] lut_7_select = {
                             in_data[46],
                             in_data[38],
                             in_data[36],
                             in_data[42],
                             in_data[6],
                             in_data[4]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [63:0] lut_8_table = 64'b0010001100000010000000000000000000111011001000110000001000000000;
    wire [5:0] lut_8_select = {
                             in_data[13],
                             in_data[29],
                             in_data[39],
                             in_data[59],
                             in_data[11],
                             in_data[23]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [63:0] lut_9_table = 64'b0000100010101111000010001000110000000000000010000000000000001000;
    wire [5:0] lut_9_select = {
                             in_data[43],
                             in_data[12],
                             in_data[49],
                             in_data[55],
                             in_data[56],
                             in_data[5]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
endmodule

